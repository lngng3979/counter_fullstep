magic
tech sky130A
magscale 1 2
timestamp 1734667522
<< checkpaint >>
rect -3932 -3932 13607 15751
<< viali >>
rect 4629 9129 4663 9163
rect 4813 8925 4847 8959
rect 5457 8925 5491 8959
rect 5273 8789 5307 8823
rect 4261 8585 4295 8619
rect 5641 8585 5675 8619
rect 4077 8517 4111 8551
rect 1593 8449 1627 8483
rect 2053 8449 2087 8483
rect 3065 8449 3099 8483
rect 4353 8449 4387 8483
rect 5549 8449 5583 8483
rect 5733 8449 5767 8483
rect 1961 8381 1995 8415
rect 2973 8381 3007 8415
rect 4445 8381 4479 8415
rect 4905 8381 4939 8415
rect 4997 8381 5031 8415
rect 5457 8381 5491 8415
rect 1409 8313 1443 8347
rect 2421 8313 2455 8347
rect 4077 8313 4111 8347
rect 4813 8313 4847 8347
rect 5273 8313 5307 8347
rect 2789 8245 2823 8279
rect 6745 8041 6779 8075
rect 4721 7973 4755 8007
rect 4261 7905 4295 7939
rect 4353 7905 4387 7939
rect 4445 7905 4479 7939
rect 4537 7905 4571 7939
rect 6009 7905 6043 7939
rect 1409 7837 1443 7871
rect 2697 7837 2731 7871
rect 2973 7837 3007 7871
rect 4905 7837 4939 7871
rect 5273 7837 5307 7871
rect 5365 7837 5399 7871
rect 5549 7837 5583 7871
rect 5917 7837 5951 7871
rect 6561 7837 6595 7871
rect 8033 7837 8067 7871
rect 2881 7769 2915 7803
rect 4997 7769 5031 7803
rect 5089 7769 5123 7803
rect 6377 7769 6411 7803
rect 1593 7701 1627 7735
rect 2513 7701 2547 7735
rect 4077 7701 4111 7735
rect 5365 7701 5399 7735
rect 6285 7701 6319 7735
rect 8217 7701 8251 7735
rect 8033 7497 8067 7531
rect 2881 7429 2915 7463
rect 5641 7361 5675 7395
rect 7205 7361 7239 7395
rect 7297 7361 7331 7395
rect 7389 7361 7423 7395
rect 7573 7361 7607 7395
rect 8217 7361 8251 7395
rect 3157 7293 3191 7327
rect 1409 7157 1443 7191
rect 4169 7157 4203 7191
rect 7021 7157 7055 7191
rect 1777 6953 1811 6987
rect 2605 6953 2639 6987
rect 4058 6953 4092 6987
rect 5549 6953 5583 6987
rect 8217 6953 8251 6987
rect 5825 6885 5859 6919
rect 3801 6817 3835 6851
rect 6469 6817 6503 6851
rect 6745 6817 6779 6851
rect 1501 6749 1535 6783
rect 2053 6749 2087 6783
rect 2421 6749 2455 6783
rect 5733 6749 5767 6783
rect 5917 6749 5951 6783
rect 6193 6749 6227 6783
rect 2237 6681 2271 6715
rect 2329 6681 2363 6715
rect 6009 6681 6043 6715
rect 6377 6613 6411 6647
rect 4905 6409 4939 6443
rect 6653 6409 6687 6443
rect 1409 6273 1443 6307
rect 1869 6273 1903 6307
rect 2513 6273 2547 6307
rect 5089 6273 5123 6307
rect 5733 6273 5767 6307
rect 6009 6273 6043 6307
rect 6193 6273 6227 6307
rect 6837 6273 6871 6307
rect 6929 6273 6963 6307
rect 7113 6273 7147 6307
rect 8033 6273 8067 6307
rect 2789 6205 2823 6239
rect 5181 6205 5215 6239
rect 5273 6205 5307 6239
rect 5365 6205 5399 6239
rect 5549 6205 5583 6239
rect 7021 6205 7055 6239
rect 1593 6137 1627 6171
rect 8217 6137 8251 6171
rect 1685 6069 1719 6103
rect 4261 6069 4295 6103
rect 2697 5865 2731 5899
rect 7665 5797 7699 5831
rect 1685 5729 1719 5763
rect 1593 5661 1627 5695
rect 2053 5661 2087 5695
rect 2201 5661 2235 5695
rect 2518 5661 2552 5695
rect 6929 5661 6963 5695
rect 7021 5661 7055 5695
rect 7297 5661 7331 5695
rect 7389 5661 7423 5695
rect 7665 5661 7699 5695
rect 8217 5661 8251 5695
rect 2329 5593 2363 5627
rect 2421 5593 2455 5627
rect 4537 5593 4571 5627
rect 7113 5593 7147 5627
rect 1961 5525 1995 5559
rect 5825 5525 5859 5559
rect 6745 5525 6779 5559
rect 8033 5525 8067 5559
rect 2237 5321 2271 5355
rect 5273 5321 5307 5355
rect 5641 5321 5675 5355
rect 8033 5321 8067 5355
rect 2053 5253 2087 5287
rect 2697 5253 2731 5287
rect 4997 5253 5031 5287
rect 7573 5253 7607 5287
rect 1409 5185 1443 5219
rect 2329 5185 2363 5219
rect 2421 5185 2455 5219
rect 3525 5185 3559 5219
rect 3709 5185 3743 5219
rect 4077 5185 4111 5219
rect 4905 5185 4939 5219
rect 5089 5185 5123 5219
rect 5181 5185 5215 5219
rect 5457 5185 5491 5219
rect 6193 5185 6227 5219
rect 6837 5185 6871 5219
rect 8217 5185 8251 5219
rect 2513 5117 2547 5151
rect 2697 5117 2731 5151
rect 5733 5117 5767 5151
rect 6561 5117 6595 5151
rect 6653 5117 6687 5151
rect 6745 5117 6779 5151
rect 1593 5049 1627 5083
rect 2053 5049 2087 5083
rect 3985 5049 4019 5083
rect 5917 5049 5951 5083
rect 7113 5049 7147 5083
rect 7297 5049 7331 5083
rect 3709 4981 3743 5015
rect 4169 4981 4203 5015
rect 6377 4981 6411 5015
rect 2329 4777 2363 4811
rect 5181 4777 5215 4811
rect 6101 4777 6135 4811
rect 6285 4777 6319 4811
rect 8217 4777 8251 4811
rect 4169 4709 4203 4743
rect 5273 4709 5307 4743
rect 2421 4641 2455 4675
rect 6469 4641 6503 4675
rect 6745 4641 6779 4675
rect 2145 4573 2179 4607
rect 2237 4573 2271 4607
rect 3801 4573 3835 4607
rect 4077 4573 4111 4607
rect 4261 4573 4295 4607
rect 4445 4573 4479 4607
rect 5733 4573 5767 4607
rect 6193 4573 6227 4607
rect 6377 4573 6411 4607
rect 5641 4505 5675 4539
rect 5917 4505 5951 4539
rect 2145 4233 2179 4267
rect 4353 4233 4387 4267
rect 3341 4165 3375 4199
rect 6377 4165 6411 4199
rect 1593 4097 1627 4131
rect 2053 4097 2087 4131
rect 3157 4097 3191 4131
rect 3525 4097 3559 4131
rect 3617 4097 3651 4131
rect 3801 4097 3835 4131
rect 4537 4097 4571 4131
rect 5181 4097 5215 4131
rect 5549 4097 5583 4131
rect 6561 4097 6595 4131
rect 6653 4097 6687 4131
rect 1685 4029 1719 4063
rect 1961 4029 1995 4063
rect 4813 4029 4847 4063
rect 4905 4029 4939 4063
rect 3709 3893 3743 3927
rect 4721 3893 4755 3927
rect 4997 3893 5031 3927
rect 5365 3893 5399 3927
rect 6377 3893 6411 3927
rect 1409 3621 1443 3655
rect 4445 3621 4479 3655
rect 2881 3553 2915 3587
rect 2973 3553 3007 3587
rect 4813 3553 4847 3587
rect 5089 3553 5123 3587
rect 1593 3485 1627 3519
rect 3065 3485 3099 3519
rect 3157 3485 3191 3519
rect 4077 3485 4111 3519
rect 4170 3485 4204 3519
rect 4721 3485 4755 3519
rect 5457 3485 5491 3519
rect 7481 3485 7515 3519
rect 2697 3349 2731 3383
rect 6745 3349 6779 3383
rect 7389 3349 7423 3383
rect 1501 3145 1535 3179
rect 8217 3145 8251 3179
rect 2973 3077 3007 3111
rect 3249 3009 3283 3043
rect 5089 3009 5123 3043
rect 5181 3009 5215 3043
rect 5365 3009 5399 3043
rect 5457 3009 5491 3043
rect 5549 3009 5583 3043
rect 5825 3009 5859 3043
rect 6009 3009 6043 3043
rect 6469 3009 6503 3043
rect 3341 2941 3375 2975
rect 4813 2941 4847 2975
rect 6745 2941 6779 2975
rect 5733 2805 5767 2839
rect 5917 2805 5951 2839
rect 3157 2601 3191 2635
rect 4997 2601 5031 2635
rect 5733 2601 5767 2635
rect 6377 2601 6411 2635
rect 7481 2601 7515 2635
rect 7849 2601 7883 2635
rect 7113 2465 7147 2499
rect 2605 2397 2639 2431
rect 2881 2397 2915 2431
rect 2973 2397 3007 2431
rect 3525 2397 3559 2431
rect 4813 2397 4847 2431
rect 5181 2397 5215 2431
rect 5457 2397 5491 2431
rect 5549 2397 5583 2431
rect 6561 2397 6595 2431
rect 6653 2397 6687 2431
rect 6929 2397 6963 2431
rect 7205 2397 7239 2431
rect 7297 2397 7331 2431
rect 7665 2397 7699 2431
rect 8217 2397 8251 2431
rect 2789 2329 2823 2363
rect 6745 2329 6779 2363
rect 3341 2261 3375 2295
rect 4629 2261 4663 2295
rect 5365 2261 5399 2295
rect 8033 2261 8067 2295
<< metal1 >>
rect 1104 9274 8556 9296
rect 1104 9222 4214 9274
rect 4266 9222 4278 9274
rect 4330 9222 4342 9274
rect 4394 9222 4406 9274
rect 4458 9222 4470 9274
rect 4522 9222 8556 9274
rect 1104 9200 8556 9222
rect 4614 9120 4620 9172
rect 4672 9120 4678 9172
rect 4798 8916 4804 8968
rect 4856 8916 4862 8968
rect 5166 8916 5172 8968
rect 5224 8956 5230 8968
rect 5445 8959 5503 8965
rect 5445 8956 5457 8959
rect 5224 8928 5457 8956
rect 5224 8916 5230 8928
rect 5445 8925 5457 8928
rect 5491 8925 5503 8959
rect 5445 8919 5503 8925
rect 5258 8780 5264 8832
rect 5316 8780 5322 8832
rect 1104 8730 8556 8752
rect 1104 8678 4874 8730
rect 4926 8678 4938 8730
rect 4990 8678 5002 8730
rect 5054 8678 5066 8730
rect 5118 8678 5130 8730
rect 5182 8678 8556 8730
rect 1104 8656 8556 8678
rect 4249 8619 4307 8625
rect 4249 8585 4261 8619
rect 4295 8616 4307 8619
rect 5626 8616 5632 8628
rect 4295 8588 5632 8616
rect 4295 8585 4307 8588
rect 4249 8579 4307 8585
rect 5626 8576 5632 8588
rect 5684 8576 5690 8628
rect 4065 8551 4123 8557
rect 2056 8520 3924 8548
rect 2056 8492 2084 8520
rect 1578 8440 1584 8492
rect 1636 8480 1642 8492
rect 1636 8452 1992 8480
rect 1636 8440 1642 8452
rect 1964 8421 1992 8452
rect 2038 8440 2044 8492
rect 2096 8440 2102 8492
rect 3053 8483 3111 8489
rect 3053 8449 3065 8483
rect 3099 8449 3111 8483
rect 3896 8480 3924 8520
rect 4065 8517 4077 8551
rect 4111 8548 4123 8551
rect 4522 8548 4528 8560
rect 4111 8520 4528 8548
rect 4111 8517 4123 8520
rect 4065 8511 4123 8517
rect 4522 8508 4528 8520
rect 4580 8548 4586 8560
rect 4580 8520 5580 8548
rect 4580 8508 4586 8520
rect 3896 8452 4200 8480
rect 3053 8443 3111 8449
rect 1949 8415 2007 8421
rect 1949 8381 1961 8415
rect 1995 8381 2007 8415
rect 2961 8415 3019 8421
rect 2961 8412 2973 8415
rect 1949 8375 2007 8381
rect 2424 8384 2973 8412
rect 1394 8304 1400 8356
rect 1452 8304 1458 8356
rect 2424 8353 2452 8384
rect 2961 8381 2973 8384
rect 3007 8381 3019 8415
rect 3068 8412 3096 8443
rect 4172 8412 4200 8452
rect 4338 8440 4344 8492
rect 4396 8440 4402 8492
rect 5552 8489 5580 8520
rect 5537 8483 5595 8489
rect 4448 8452 5304 8480
rect 4448 8421 4476 8452
rect 4433 8415 4491 8421
rect 4433 8412 4445 8415
rect 3068 8384 4108 8412
rect 4172 8384 4445 8412
rect 2961 8375 3019 8381
rect 4080 8353 4108 8384
rect 4433 8381 4445 8384
rect 4479 8381 4491 8415
rect 4433 8375 4491 8381
rect 4522 8372 4528 8424
rect 4580 8412 4586 8424
rect 4893 8415 4951 8421
rect 4893 8412 4905 8415
rect 4580 8384 4905 8412
rect 4580 8372 4586 8384
rect 4893 8381 4905 8384
rect 4939 8381 4951 8415
rect 4893 8375 4951 8381
rect 4982 8372 4988 8424
rect 5040 8372 5046 8424
rect 2409 8347 2467 8353
rect 2409 8313 2421 8347
rect 2455 8313 2467 8347
rect 2409 8307 2467 8313
rect 4065 8347 4123 8353
rect 4065 8313 4077 8347
rect 4111 8313 4123 8347
rect 4065 8307 4123 8313
rect 4801 8347 4859 8353
rect 4801 8313 4813 8347
rect 4847 8344 4859 8347
rect 5000 8344 5028 8372
rect 5276 8353 5304 8452
rect 5537 8449 5549 8483
rect 5583 8449 5595 8483
rect 5537 8443 5595 8449
rect 5721 8483 5779 8489
rect 5721 8449 5733 8483
rect 5767 8449 5779 8483
rect 5721 8443 5779 8449
rect 5445 8415 5503 8421
rect 5445 8381 5457 8415
rect 5491 8412 5503 8415
rect 5736 8412 5764 8443
rect 5491 8384 5764 8412
rect 5491 8381 5503 8384
rect 5445 8375 5503 8381
rect 4847 8316 5028 8344
rect 5261 8347 5319 8353
rect 4847 8313 4859 8316
rect 4801 8307 4859 8313
rect 5261 8313 5273 8347
rect 5307 8344 5319 8347
rect 5902 8344 5908 8356
rect 5307 8316 5908 8344
rect 5307 8313 5319 8316
rect 5261 8307 5319 8313
rect 5902 8304 5908 8316
rect 5960 8304 5966 8356
rect 2774 8236 2780 8288
rect 2832 8236 2838 8288
rect 4338 8236 4344 8288
rect 4396 8276 4402 8288
rect 5442 8276 5448 8288
rect 4396 8248 5448 8276
rect 4396 8236 4402 8248
rect 5442 8236 5448 8248
rect 5500 8236 5506 8288
rect 1104 8186 8556 8208
rect 1104 8134 4214 8186
rect 4266 8134 4278 8186
rect 4330 8134 4342 8186
rect 4394 8134 4406 8186
rect 4458 8134 4470 8186
rect 4522 8134 8556 8186
rect 1104 8112 8556 8134
rect 6733 8075 6791 8081
rect 6733 8072 6745 8075
rect 4264 8044 6745 8072
rect 4264 7945 4292 8044
rect 6733 8041 6745 8044
rect 6779 8041 6791 8075
rect 6733 8035 6791 8041
rect 4709 8007 4767 8013
rect 4709 8004 4721 8007
rect 4540 7976 4721 8004
rect 4249 7939 4307 7945
rect 4249 7905 4261 7939
rect 4295 7905 4307 7939
rect 4249 7899 4307 7905
rect 4338 7896 4344 7948
rect 4396 7896 4402 7948
rect 4430 7896 4436 7948
rect 4488 7896 4494 7948
rect 4540 7945 4568 7976
rect 4709 7973 4721 7976
rect 4755 7973 4767 8007
rect 5258 8004 5264 8016
rect 4709 7967 4767 7973
rect 4908 7976 5264 8004
rect 4525 7939 4583 7945
rect 4525 7905 4537 7939
rect 4571 7905 4583 7939
rect 4525 7899 4583 7905
rect 842 7828 848 7880
rect 900 7868 906 7880
rect 1397 7871 1455 7877
rect 1397 7868 1409 7871
rect 900 7840 1409 7868
rect 900 7828 906 7840
rect 1397 7837 1409 7840
rect 1443 7837 1455 7871
rect 1397 7831 1455 7837
rect 2682 7828 2688 7880
rect 2740 7828 2746 7880
rect 2774 7828 2780 7880
rect 2832 7868 2838 7880
rect 4908 7877 4936 7976
rect 5258 7964 5264 7976
rect 5316 7964 5322 8016
rect 5644 7976 6592 8004
rect 5644 7948 5672 7976
rect 4982 7896 4988 7948
rect 5040 7936 5046 7948
rect 5626 7936 5632 7948
rect 5040 7908 5304 7936
rect 5040 7896 5046 7908
rect 2961 7871 3019 7877
rect 2961 7868 2973 7871
rect 2832 7840 2973 7868
rect 2832 7828 2838 7840
rect 2961 7837 2973 7840
rect 3007 7837 3019 7871
rect 2961 7831 3019 7837
rect 4893 7871 4951 7877
rect 4893 7837 4905 7871
rect 4939 7837 4951 7871
rect 4893 7831 4951 7837
rect 5166 7828 5172 7880
rect 5224 7828 5230 7880
rect 5276 7877 5304 7908
rect 5368 7908 5632 7936
rect 5368 7877 5396 7908
rect 5626 7896 5632 7908
rect 5684 7896 5690 7948
rect 5994 7896 6000 7948
rect 6052 7896 6058 7948
rect 5261 7871 5319 7877
rect 5261 7837 5273 7871
rect 5307 7837 5319 7871
rect 5261 7831 5319 7837
rect 5353 7871 5411 7877
rect 5353 7837 5365 7871
rect 5399 7837 5411 7871
rect 5353 7831 5411 7837
rect 2590 7760 2596 7812
rect 2648 7800 2654 7812
rect 2869 7803 2927 7809
rect 2869 7800 2881 7803
rect 2648 7772 2881 7800
rect 2648 7760 2654 7772
rect 2869 7769 2881 7772
rect 2915 7800 2927 7803
rect 4430 7800 4436 7812
rect 2915 7772 4436 7800
rect 2915 7769 2927 7772
rect 2869 7763 2927 7769
rect 4430 7760 4436 7772
rect 4488 7760 4494 7812
rect 4798 7760 4804 7812
rect 4856 7800 4862 7812
rect 4985 7803 5043 7809
rect 4985 7800 4997 7803
rect 4856 7772 4997 7800
rect 4856 7760 4862 7772
rect 4985 7769 4997 7772
rect 5031 7769 5043 7803
rect 4985 7763 5043 7769
rect 5077 7803 5135 7809
rect 5077 7769 5089 7803
rect 5123 7800 5135 7803
rect 5184 7800 5212 7828
rect 5123 7772 5212 7800
rect 5276 7800 5304 7831
rect 5442 7828 5448 7880
rect 5500 7868 5506 7880
rect 5537 7871 5595 7877
rect 5537 7868 5549 7871
rect 5500 7840 5549 7868
rect 5500 7828 5506 7840
rect 5537 7837 5549 7840
rect 5583 7868 5595 7871
rect 5583 7840 5764 7868
rect 5583 7837 5595 7840
rect 5537 7831 5595 7837
rect 5626 7800 5632 7812
rect 5276 7772 5632 7800
rect 5123 7769 5135 7772
rect 5077 7763 5135 7769
rect 5626 7760 5632 7772
rect 5684 7760 5690 7812
rect 1581 7735 1639 7741
rect 1581 7701 1593 7735
rect 1627 7732 1639 7735
rect 2406 7732 2412 7744
rect 1627 7704 2412 7732
rect 1627 7701 1639 7704
rect 1581 7695 1639 7701
rect 2406 7692 2412 7704
rect 2464 7692 2470 7744
rect 2501 7735 2559 7741
rect 2501 7701 2513 7735
rect 2547 7732 2559 7735
rect 2774 7732 2780 7744
rect 2547 7704 2780 7732
rect 2547 7701 2559 7704
rect 2501 7695 2559 7701
rect 2774 7692 2780 7704
rect 2832 7692 2838 7744
rect 3878 7692 3884 7744
rect 3936 7732 3942 7744
rect 4065 7735 4123 7741
rect 4065 7732 4077 7735
rect 3936 7704 4077 7732
rect 3936 7692 3942 7704
rect 4065 7701 4077 7704
rect 4111 7701 4123 7735
rect 4065 7695 4123 7701
rect 4338 7692 4344 7744
rect 4396 7732 4402 7744
rect 5353 7735 5411 7741
rect 5353 7732 5365 7735
rect 4396 7704 5365 7732
rect 4396 7692 4402 7704
rect 5353 7701 5365 7704
rect 5399 7701 5411 7735
rect 5736 7732 5764 7840
rect 5902 7828 5908 7880
rect 5960 7828 5966 7880
rect 6564 7877 6592 7976
rect 6549 7871 6607 7877
rect 6549 7837 6561 7871
rect 6595 7837 6607 7871
rect 6549 7831 6607 7837
rect 6822 7828 6828 7880
rect 6880 7868 6886 7880
rect 8021 7871 8079 7877
rect 8021 7868 8033 7871
rect 6880 7840 8033 7868
rect 6880 7828 6886 7840
rect 8021 7837 8033 7840
rect 8067 7837 8079 7871
rect 8021 7831 8079 7837
rect 6365 7803 6423 7809
rect 6365 7800 6377 7803
rect 6104 7772 6377 7800
rect 6104 7732 6132 7772
rect 6365 7769 6377 7772
rect 6411 7769 6423 7803
rect 6365 7763 6423 7769
rect 5736 7704 6132 7732
rect 5353 7695 5411 7701
rect 6270 7692 6276 7744
rect 6328 7692 6334 7744
rect 8202 7692 8208 7744
rect 8260 7692 8266 7744
rect 1104 7642 8556 7664
rect 1104 7590 4874 7642
rect 4926 7590 4938 7642
rect 4990 7590 5002 7642
rect 5054 7590 5066 7642
rect 5118 7590 5130 7642
rect 5182 7590 8556 7642
rect 1104 7568 8556 7590
rect 3234 7528 3240 7540
rect 2700 7500 3240 7528
rect 2700 7460 2728 7500
rect 3234 7488 3240 7500
rect 3292 7488 3298 7540
rect 4798 7488 4804 7540
rect 4856 7528 4862 7540
rect 7282 7528 7288 7540
rect 4856 7500 7288 7528
rect 4856 7488 4862 7500
rect 7282 7488 7288 7500
rect 7340 7488 7346 7540
rect 8021 7531 8079 7537
rect 8021 7497 8033 7531
rect 8067 7497 8079 7531
rect 8021 7491 8079 7497
rect 2438 7432 2728 7460
rect 2774 7420 2780 7472
rect 2832 7460 2838 7472
rect 2869 7463 2927 7469
rect 2869 7460 2881 7463
rect 2832 7432 2881 7460
rect 2832 7420 2838 7432
rect 2869 7429 2881 7432
rect 2915 7429 2927 7463
rect 8036 7460 8064 7491
rect 2869 7423 2927 7429
rect 7208 7432 8064 7460
rect 5629 7395 5687 7401
rect 5629 7361 5641 7395
rect 5675 7392 5687 7395
rect 5810 7392 5816 7404
rect 5675 7364 5816 7392
rect 5675 7361 5687 7364
rect 5629 7355 5687 7361
rect 5810 7352 5816 7364
rect 5868 7352 5874 7404
rect 7208 7401 7236 7432
rect 7193 7395 7251 7401
rect 7193 7361 7205 7395
rect 7239 7361 7251 7395
rect 7193 7355 7251 7361
rect 7282 7352 7288 7404
rect 7340 7352 7346 7404
rect 7377 7395 7435 7401
rect 7377 7361 7389 7395
rect 7423 7392 7435 7395
rect 7466 7392 7472 7404
rect 7423 7364 7472 7392
rect 7423 7361 7435 7364
rect 7377 7355 7435 7361
rect 7466 7352 7472 7364
rect 7524 7352 7530 7404
rect 7561 7395 7619 7401
rect 7561 7361 7573 7395
rect 7607 7361 7619 7395
rect 7561 7355 7619 7361
rect 3142 7284 3148 7336
rect 3200 7324 3206 7336
rect 3200 7296 4108 7324
rect 3200 7284 3206 7296
rect 4080 7200 4108 7296
rect 5994 7284 6000 7336
rect 6052 7324 6058 7336
rect 6822 7324 6828 7336
rect 6052 7296 6828 7324
rect 6052 7284 6058 7296
rect 6822 7284 6828 7296
rect 6880 7324 6886 7336
rect 7576 7324 7604 7355
rect 8202 7352 8208 7404
rect 8260 7352 8266 7404
rect 6880 7296 7604 7324
rect 6880 7284 6886 7296
rect 5258 7216 5264 7268
rect 5316 7256 5322 7268
rect 7466 7256 7472 7268
rect 5316 7228 7472 7256
rect 5316 7216 5322 7228
rect 7466 7216 7472 7228
rect 7524 7216 7530 7268
rect 1397 7191 1455 7197
rect 1397 7157 1409 7191
rect 1443 7188 1455 7191
rect 1578 7188 1584 7200
rect 1443 7160 1584 7188
rect 1443 7157 1455 7160
rect 1397 7151 1455 7157
rect 1578 7148 1584 7160
rect 1636 7148 1642 7200
rect 4062 7148 4068 7200
rect 4120 7188 4126 7200
rect 4157 7191 4215 7197
rect 4157 7188 4169 7191
rect 4120 7160 4169 7188
rect 4120 7148 4126 7160
rect 4157 7157 4169 7160
rect 4203 7157 4215 7191
rect 4157 7151 4215 7157
rect 7009 7191 7067 7197
rect 7009 7157 7021 7191
rect 7055 7188 7067 7191
rect 7098 7188 7104 7200
rect 7055 7160 7104 7188
rect 7055 7157 7067 7160
rect 7009 7151 7067 7157
rect 7098 7148 7104 7160
rect 7156 7148 7162 7200
rect 1104 7098 8556 7120
rect 1104 7046 4214 7098
rect 4266 7046 4278 7098
rect 4330 7046 4342 7098
rect 4394 7046 4406 7098
rect 4458 7046 4470 7098
rect 4522 7046 8556 7098
rect 1104 7024 8556 7046
rect 1762 6944 1768 6996
rect 1820 6984 1826 6996
rect 2038 6984 2044 6996
rect 1820 6956 2044 6984
rect 1820 6944 1826 6956
rect 2038 6944 2044 6956
rect 2096 6944 2102 6996
rect 2593 6987 2651 6993
rect 2593 6953 2605 6987
rect 2639 6984 2651 6987
rect 2682 6984 2688 6996
rect 2639 6956 2688 6984
rect 2639 6953 2651 6956
rect 2593 6947 2651 6953
rect 2682 6944 2688 6956
rect 2740 6944 2746 6996
rect 3878 6944 3884 6996
rect 3936 6984 3942 6996
rect 4046 6987 4104 6993
rect 4046 6984 4058 6987
rect 3936 6956 4058 6984
rect 3936 6944 3942 6956
rect 4046 6953 4058 6956
rect 4092 6953 4104 6987
rect 4046 6947 4104 6953
rect 5537 6987 5595 6993
rect 5537 6953 5549 6987
rect 5583 6984 5595 6987
rect 5626 6984 5632 6996
rect 5583 6956 5632 6984
rect 5583 6953 5595 6956
rect 5537 6947 5595 6953
rect 5626 6944 5632 6956
rect 5684 6944 5690 6996
rect 6822 6944 6828 6996
rect 6880 6984 6886 6996
rect 8205 6987 8263 6993
rect 8205 6984 8217 6987
rect 6880 6956 8217 6984
rect 6880 6944 6886 6956
rect 8205 6953 8217 6956
rect 8251 6953 8263 6987
rect 8205 6947 8263 6953
rect 5813 6919 5871 6925
rect 5813 6885 5825 6919
rect 5859 6916 5871 6919
rect 5902 6916 5908 6928
rect 5859 6888 5908 6916
rect 5859 6885 5871 6888
rect 5813 6879 5871 6885
rect 5902 6876 5908 6888
rect 5960 6876 5966 6928
rect 3789 6851 3847 6857
rect 3789 6817 3801 6851
rect 3835 6848 3847 6851
rect 4062 6848 4068 6860
rect 3835 6820 4068 6848
rect 3835 6817 3847 6820
rect 3789 6811 3847 6817
rect 4062 6808 4068 6820
rect 4120 6848 4126 6860
rect 6457 6851 6515 6857
rect 6457 6848 6469 6851
rect 4120 6820 6469 6848
rect 4120 6808 4126 6820
rect 6457 6817 6469 6820
rect 6503 6817 6515 6851
rect 6457 6811 6515 6817
rect 6730 6808 6736 6860
rect 6788 6808 6794 6860
rect 934 6740 940 6792
rect 992 6780 998 6792
rect 1489 6783 1547 6789
rect 1489 6780 1501 6783
rect 992 6752 1501 6780
rect 992 6740 998 6752
rect 1489 6749 1501 6752
rect 1535 6749 1547 6783
rect 1489 6743 1547 6749
rect 1578 6740 1584 6792
rect 1636 6780 1642 6792
rect 2041 6783 2099 6789
rect 2041 6780 2053 6783
rect 1636 6752 2053 6780
rect 1636 6740 1642 6752
rect 2041 6749 2053 6752
rect 2087 6749 2099 6783
rect 2041 6743 2099 6749
rect 2406 6740 2412 6792
rect 2464 6740 2470 6792
rect 5718 6740 5724 6792
rect 5776 6740 5782 6792
rect 5905 6783 5963 6789
rect 5905 6749 5917 6783
rect 5951 6780 5963 6783
rect 6181 6783 6239 6789
rect 6181 6780 6193 6783
rect 5951 6752 6193 6780
rect 5951 6749 5963 6752
rect 5905 6743 5963 6749
rect 6181 6749 6193 6752
rect 6227 6780 6239 6783
rect 6270 6780 6276 6792
rect 6227 6752 6276 6780
rect 6227 6749 6239 6752
rect 6181 6743 6239 6749
rect 6270 6740 6276 6752
rect 6328 6740 6334 6792
rect 2222 6672 2228 6724
rect 2280 6672 2286 6724
rect 2317 6715 2375 6721
rect 2317 6681 2329 6715
rect 2363 6712 2375 6715
rect 2363 6684 2452 6712
rect 2363 6681 2375 6684
rect 2317 6675 2375 6681
rect 2424 6656 2452 6684
rect 3234 6672 3240 6724
rect 3292 6712 3298 6724
rect 5736 6712 5764 6740
rect 5997 6715 6055 6721
rect 5997 6712 6009 6715
rect 3292 6684 4554 6712
rect 5736 6684 6009 6712
rect 3292 6672 3298 6684
rect 2406 6604 2412 6656
rect 2464 6604 2470 6656
rect 4448 6644 4476 6684
rect 5997 6681 6009 6684
rect 6043 6681 6055 6715
rect 5997 6675 6055 6681
rect 6104 6684 7222 6712
rect 6104 6644 6132 6684
rect 4448 6616 6132 6644
rect 6365 6647 6423 6653
rect 6365 6613 6377 6647
rect 6411 6644 6423 6647
rect 6822 6644 6828 6656
rect 6411 6616 6828 6644
rect 6411 6613 6423 6616
rect 6365 6607 6423 6613
rect 6822 6604 6828 6616
rect 6880 6604 6886 6656
rect 7116 6644 7144 6684
rect 7374 6644 7380 6656
rect 7116 6616 7380 6644
rect 7374 6604 7380 6616
rect 7432 6604 7438 6656
rect 1104 6554 8556 6576
rect 1104 6502 4874 6554
rect 4926 6502 4938 6554
rect 4990 6502 5002 6554
rect 5054 6502 5066 6554
rect 5118 6502 5130 6554
rect 5182 6502 8556 6554
rect 1104 6480 8556 6502
rect 3142 6440 3148 6452
rect 2516 6412 3148 6440
rect 842 6264 848 6316
rect 900 6304 906 6316
rect 1397 6307 1455 6313
rect 1397 6304 1409 6307
rect 900 6276 1409 6304
rect 900 6264 906 6276
rect 1397 6273 1409 6276
rect 1443 6273 1455 6307
rect 1397 6267 1455 6273
rect 1854 6264 1860 6316
rect 1912 6264 1918 6316
rect 2516 6313 2544 6412
rect 3142 6400 3148 6412
rect 3200 6400 3206 6452
rect 4893 6443 4951 6449
rect 4893 6409 4905 6443
rect 4939 6440 4951 6443
rect 5350 6440 5356 6452
rect 4939 6412 5356 6440
rect 4939 6409 4951 6412
rect 4893 6403 4951 6409
rect 5350 6400 5356 6412
rect 5408 6400 5414 6452
rect 6270 6440 6276 6452
rect 5644 6412 6276 6440
rect 3234 6332 3240 6384
rect 3292 6332 3298 6384
rect 2501 6307 2559 6313
rect 2501 6273 2513 6307
rect 2547 6273 2559 6307
rect 2501 6267 2559 6273
rect 5077 6307 5135 6313
rect 5077 6273 5089 6307
rect 5123 6304 5135 6307
rect 5644 6304 5672 6412
rect 6270 6400 6276 6412
rect 6328 6400 6334 6452
rect 6641 6443 6699 6449
rect 6641 6409 6653 6443
rect 6687 6440 6699 6443
rect 6730 6440 6736 6452
rect 6687 6412 6736 6440
rect 6687 6409 6699 6412
rect 6641 6403 6699 6409
rect 6730 6400 6736 6412
rect 6788 6400 6794 6452
rect 5902 6332 5908 6384
rect 5960 6372 5966 6384
rect 5960 6344 6960 6372
rect 5960 6332 5966 6344
rect 5123 6276 5672 6304
rect 5721 6307 5779 6313
rect 5123 6273 5135 6276
rect 5077 6267 5135 6273
rect 5721 6273 5733 6307
rect 5767 6273 5779 6307
rect 5721 6267 5779 6273
rect 2774 6196 2780 6248
rect 2832 6196 2838 6248
rect 5166 6196 5172 6248
rect 5224 6196 5230 6248
rect 5258 6196 5264 6248
rect 5316 6196 5322 6248
rect 5353 6239 5411 6245
rect 5353 6205 5365 6239
rect 5399 6236 5411 6239
rect 5537 6239 5595 6245
rect 5537 6236 5549 6239
rect 5399 6208 5549 6236
rect 5399 6205 5411 6208
rect 5353 6199 5411 6205
rect 5537 6205 5549 6208
rect 5583 6205 5595 6239
rect 5537 6199 5595 6205
rect 5626 6196 5632 6248
rect 5684 6236 5690 6248
rect 5736 6236 5764 6267
rect 5994 6264 6000 6316
rect 6052 6264 6058 6316
rect 6178 6264 6184 6316
rect 6236 6264 6242 6316
rect 6822 6264 6828 6316
rect 6880 6264 6886 6316
rect 6932 6313 6960 6344
rect 6917 6307 6975 6313
rect 6917 6273 6929 6307
rect 6963 6273 6975 6307
rect 6917 6267 6975 6273
rect 7098 6264 7104 6316
rect 7156 6264 7162 6316
rect 8018 6264 8024 6316
rect 8076 6264 8082 6316
rect 5684 6208 5764 6236
rect 5684 6196 5690 6208
rect 6730 6196 6736 6248
rect 6788 6236 6794 6248
rect 7009 6239 7067 6245
rect 7009 6236 7021 6239
rect 6788 6208 7021 6236
rect 6788 6196 6794 6208
rect 7009 6205 7021 6208
rect 7055 6205 7067 6239
rect 7009 6199 7067 6205
rect 1581 6171 1639 6177
rect 1581 6137 1593 6171
rect 1627 6168 1639 6171
rect 2498 6168 2504 6180
rect 1627 6140 2504 6168
rect 1627 6137 1639 6140
rect 1581 6131 1639 6137
rect 2498 6128 2504 6140
rect 2556 6128 2562 6180
rect 8202 6128 8208 6180
rect 8260 6128 8266 6180
rect 1670 6060 1676 6112
rect 1728 6060 1734 6112
rect 3786 6060 3792 6112
rect 3844 6100 3850 6112
rect 4249 6103 4307 6109
rect 4249 6100 4261 6103
rect 3844 6072 4261 6100
rect 3844 6060 3850 6072
rect 4249 6069 4261 6072
rect 4295 6069 4307 6103
rect 4249 6063 4307 6069
rect 1104 6010 8556 6032
rect 1104 5958 4214 6010
rect 4266 5958 4278 6010
rect 4330 5958 4342 6010
rect 4394 5958 4406 6010
rect 4458 5958 4470 6010
rect 4522 5958 8556 6010
rect 1104 5936 8556 5958
rect 2685 5899 2743 5905
rect 2685 5865 2697 5899
rect 2731 5896 2743 5899
rect 2774 5896 2780 5908
rect 2731 5868 2780 5896
rect 2731 5865 2743 5868
rect 2685 5859 2743 5865
rect 2774 5856 2780 5868
rect 2832 5856 2838 5908
rect 7466 5788 7472 5840
rect 7524 5828 7530 5840
rect 7653 5831 7711 5837
rect 7653 5828 7665 5831
rect 7524 5800 7665 5828
rect 7524 5788 7530 5800
rect 7653 5797 7665 5800
rect 7699 5797 7711 5831
rect 7653 5791 7711 5797
rect 1673 5763 1731 5769
rect 1673 5729 1685 5763
rect 1719 5760 1731 5763
rect 1854 5760 1860 5772
rect 1719 5732 1860 5760
rect 1719 5729 1731 5732
rect 1673 5723 1731 5729
rect 1854 5720 1860 5732
rect 1912 5760 1918 5772
rect 3786 5760 3792 5772
rect 1912 5732 3792 5760
rect 1912 5720 1918 5732
rect 1581 5695 1639 5701
rect 1581 5661 1593 5695
rect 1627 5692 1639 5695
rect 1762 5692 1768 5704
rect 1627 5664 1768 5692
rect 1627 5661 1639 5664
rect 1581 5655 1639 5661
rect 1762 5652 1768 5664
rect 1820 5652 1826 5704
rect 2038 5652 2044 5704
rect 2096 5652 2102 5704
rect 2240 5701 2268 5732
rect 3786 5720 3792 5732
rect 3844 5720 3850 5772
rect 6178 5720 6184 5772
rect 6236 5760 6242 5772
rect 8018 5760 8024 5772
rect 6236 5732 8024 5760
rect 6236 5720 6242 5732
rect 2189 5695 2268 5701
rect 2189 5661 2201 5695
rect 2235 5664 2268 5695
rect 2235 5661 2247 5664
rect 2189 5655 2247 5661
rect 2498 5652 2504 5704
rect 2556 5701 2562 5704
rect 2556 5692 2564 5701
rect 2556 5664 2601 5692
rect 2556 5655 2564 5664
rect 2556 5652 2562 5655
rect 6914 5652 6920 5704
rect 6972 5652 6978 5704
rect 7009 5695 7067 5701
rect 7009 5661 7021 5695
rect 7055 5692 7067 5695
rect 7190 5692 7196 5704
rect 7055 5664 7196 5692
rect 7055 5661 7067 5664
rect 7009 5655 7067 5661
rect 7190 5652 7196 5664
rect 7248 5652 7254 5704
rect 7300 5701 7328 5732
rect 8018 5720 8024 5732
rect 8076 5720 8082 5772
rect 7285 5695 7343 5701
rect 7285 5661 7297 5695
rect 7331 5661 7343 5695
rect 7285 5655 7343 5661
rect 7377 5695 7435 5701
rect 7377 5661 7389 5695
rect 7423 5661 7435 5695
rect 7377 5655 7435 5661
rect 2317 5627 2375 5633
rect 2317 5593 2329 5627
rect 2363 5593 2375 5627
rect 2317 5587 2375 5593
rect 1946 5516 1952 5568
rect 2004 5516 2010 5568
rect 2222 5516 2228 5568
rect 2280 5556 2286 5568
rect 2332 5556 2360 5587
rect 2406 5584 2412 5636
rect 2464 5624 2470 5636
rect 3234 5624 3240 5636
rect 2464 5596 3240 5624
rect 2464 5584 2470 5596
rect 3234 5584 3240 5596
rect 3292 5584 3298 5636
rect 4525 5627 4583 5633
rect 4525 5593 4537 5627
rect 4571 5624 4583 5627
rect 4614 5624 4620 5636
rect 4571 5596 4620 5624
rect 4571 5593 4583 5596
rect 4525 5587 4583 5593
rect 4614 5584 4620 5596
rect 4672 5584 4678 5636
rect 7101 5627 7159 5633
rect 7101 5593 7113 5627
rect 7147 5593 7159 5627
rect 7208 5624 7236 5652
rect 7392 5624 7420 5655
rect 7650 5652 7656 5704
rect 7708 5692 7714 5704
rect 7708 5664 8064 5692
rect 7708 5652 7714 5664
rect 7208 5596 7420 5624
rect 7101 5587 7159 5593
rect 5074 5556 5080 5568
rect 2280 5528 5080 5556
rect 2280 5516 2286 5528
rect 5074 5516 5080 5528
rect 5132 5556 5138 5568
rect 5442 5556 5448 5568
rect 5132 5528 5448 5556
rect 5132 5516 5138 5528
rect 5442 5516 5448 5528
rect 5500 5516 5506 5568
rect 5810 5516 5816 5568
rect 5868 5516 5874 5568
rect 6733 5559 6791 5565
rect 6733 5525 6745 5559
rect 6779 5556 6791 5559
rect 6822 5556 6828 5568
rect 6779 5528 6828 5556
rect 6779 5525 6791 5528
rect 6733 5519 6791 5525
rect 6822 5516 6828 5528
rect 6880 5516 6886 5568
rect 7116 5556 7144 5587
rect 7466 5556 7472 5568
rect 7116 5528 7472 5556
rect 7466 5516 7472 5528
rect 7524 5516 7530 5568
rect 8036 5565 8064 5664
rect 8202 5652 8208 5704
rect 8260 5652 8266 5704
rect 8021 5559 8079 5565
rect 8021 5525 8033 5559
rect 8067 5525 8079 5559
rect 8021 5519 8079 5525
rect 1104 5466 8556 5488
rect 1104 5414 4874 5466
rect 4926 5414 4938 5466
rect 4990 5414 5002 5466
rect 5054 5414 5066 5466
rect 5118 5414 5130 5466
rect 5182 5414 8556 5466
rect 1104 5392 8556 5414
rect 1946 5312 1952 5364
rect 2004 5352 2010 5364
rect 2225 5355 2283 5361
rect 2225 5352 2237 5355
rect 2004 5324 2237 5352
rect 2004 5312 2010 5324
rect 2225 5321 2237 5324
rect 2271 5352 2283 5355
rect 2271 5324 2820 5352
rect 2271 5321 2283 5324
rect 2225 5315 2283 5321
rect 2041 5287 2099 5293
rect 2041 5253 2053 5287
rect 2087 5284 2099 5287
rect 2685 5287 2743 5293
rect 2685 5284 2697 5287
rect 2087 5256 2697 5284
rect 2087 5253 2099 5256
rect 2041 5247 2099 5253
rect 2685 5253 2697 5256
rect 2731 5253 2743 5287
rect 2685 5247 2743 5253
rect 842 5176 848 5228
rect 900 5216 906 5228
rect 1397 5219 1455 5225
rect 1397 5216 1409 5219
rect 900 5188 1409 5216
rect 900 5176 906 5188
rect 1397 5185 1409 5188
rect 1443 5185 1455 5219
rect 1397 5179 1455 5185
rect 2314 5176 2320 5228
rect 2372 5176 2378 5228
rect 2409 5219 2467 5225
rect 2409 5185 2421 5219
rect 2455 5216 2467 5219
rect 2792 5216 2820 5324
rect 4890 5312 4896 5364
rect 4948 5352 4954 5364
rect 5261 5355 5319 5361
rect 5261 5352 5273 5355
rect 4948 5324 5273 5352
rect 4948 5312 4954 5324
rect 5261 5321 5273 5324
rect 5307 5352 5319 5355
rect 5350 5352 5356 5364
rect 5307 5324 5356 5352
rect 5307 5321 5319 5324
rect 5261 5315 5319 5321
rect 5350 5312 5356 5324
rect 5408 5312 5414 5364
rect 5629 5355 5687 5361
rect 5629 5321 5641 5355
rect 5675 5352 5687 5355
rect 5718 5352 5724 5364
rect 5675 5324 5724 5352
rect 5675 5321 5687 5324
rect 5629 5315 5687 5321
rect 5718 5312 5724 5324
rect 5776 5312 5782 5364
rect 6914 5312 6920 5364
rect 6972 5352 6978 5364
rect 8021 5355 8079 5361
rect 8021 5352 8033 5355
rect 6972 5324 8033 5352
rect 6972 5312 6978 5324
rect 8021 5321 8033 5324
rect 8067 5321 8079 5355
rect 8021 5315 8079 5321
rect 4985 5287 5043 5293
rect 3160 5256 4108 5284
rect 3160 5216 3188 5256
rect 2455 5188 3188 5216
rect 3513 5219 3571 5225
rect 2455 5185 2467 5188
rect 2409 5179 2467 5185
rect 3513 5185 3525 5219
rect 3559 5185 3571 5219
rect 3513 5179 3571 5185
rect 3697 5219 3755 5225
rect 3697 5185 3709 5219
rect 3743 5216 3755 5219
rect 3786 5216 3792 5228
rect 3743 5188 3792 5216
rect 3743 5185 3755 5188
rect 3697 5179 3755 5185
rect 2332 5148 2360 5176
rect 2501 5151 2559 5157
rect 2501 5148 2513 5151
rect 1596 5120 2268 5148
rect 2332 5120 2513 5148
rect 1596 5089 1624 5120
rect 1581 5083 1639 5089
rect 1581 5049 1593 5083
rect 1627 5049 1639 5083
rect 1581 5043 1639 5049
rect 2038 5040 2044 5092
rect 2096 5040 2102 5092
rect 2240 5080 2268 5120
rect 2501 5117 2513 5120
rect 2547 5117 2559 5151
rect 2501 5111 2559 5117
rect 2590 5108 2596 5160
rect 2648 5148 2654 5160
rect 2685 5151 2743 5157
rect 2685 5148 2697 5151
rect 2648 5120 2697 5148
rect 2648 5108 2654 5120
rect 2685 5117 2697 5120
rect 2731 5117 2743 5151
rect 2685 5111 2743 5117
rect 2774 5108 2780 5160
rect 2832 5148 2838 5160
rect 3528 5148 3556 5179
rect 3786 5176 3792 5188
rect 3844 5176 3850 5228
rect 4080 5225 4108 5256
rect 4985 5253 4997 5287
rect 5031 5284 5043 5287
rect 5031 5256 5212 5284
rect 5031 5253 5043 5256
rect 4985 5247 5043 5253
rect 5184 5228 5212 5256
rect 7282 5244 7288 5296
rect 7340 5284 7346 5296
rect 7561 5287 7619 5293
rect 7561 5284 7573 5287
rect 7340 5256 7573 5284
rect 7340 5244 7346 5256
rect 7561 5253 7573 5256
rect 7607 5253 7619 5287
rect 7561 5247 7619 5253
rect 4065 5219 4123 5225
rect 4065 5185 4077 5219
rect 4111 5185 4123 5219
rect 4065 5179 4123 5185
rect 4893 5219 4951 5225
rect 4893 5185 4905 5219
rect 4939 5185 4951 5219
rect 4893 5179 4951 5185
rect 2832 5120 3556 5148
rect 4908 5148 4936 5179
rect 5074 5176 5080 5228
rect 5132 5176 5138 5228
rect 5166 5176 5172 5228
rect 5224 5176 5230 5228
rect 5445 5219 5503 5225
rect 5445 5185 5457 5219
rect 5491 5185 5503 5219
rect 5445 5179 5503 5185
rect 5460 5148 5488 5179
rect 5626 5176 5632 5228
rect 5684 5216 5690 5228
rect 6181 5219 6239 5225
rect 6181 5216 6193 5219
rect 5684 5188 6193 5216
rect 5684 5176 5690 5188
rect 6181 5185 6193 5188
rect 6227 5185 6239 5219
rect 6181 5179 6239 5185
rect 6822 5176 6828 5228
rect 6880 5176 6886 5228
rect 6914 5176 6920 5228
rect 6972 5216 6978 5228
rect 7300 5216 7328 5244
rect 6972 5188 7328 5216
rect 6972 5176 6978 5188
rect 8202 5176 8208 5228
rect 8260 5176 8266 5228
rect 5721 5151 5779 5157
rect 5721 5148 5733 5151
rect 4908 5120 5733 5148
rect 2832 5108 2838 5120
rect 5721 5117 5733 5120
rect 5767 5117 5779 5151
rect 5721 5111 5779 5117
rect 6270 5108 6276 5160
rect 6328 5148 6334 5160
rect 6549 5151 6607 5157
rect 6549 5148 6561 5151
rect 6328 5120 6561 5148
rect 6328 5108 6334 5120
rect 6549 5117 6561 5120
rect 6595 5117 6607 5151
rect 6549 5111 6607 5117
rect 6641 5151 6699 5157
rect 6641 5117 6653 5151
rect 6687 5117 6699 5151
rect 6641 5111 6699 5117
rect 2406 5080 2412 5092
rect 2240 5052 2412 5080
rect 2406 5040 2412 5052
rect 2464 5040 2470 5092
rect 3878 5080 3884 5092
rect 3620 5052 3884 5080
rect 1762 4972 1768 5024
rect 1820 5012 1826 5024
rect 3620 5012 3648 5052
rect 3878 5040 3884 5052
rect 3936 5080 3942 5092
rect 3973 5083 4031 5089
rect 3973 5080 3985 5083
rect 3936 5052 3985 5080
rect 3936 5040 3942 5052
rect 3973 5049 3985 5052
rect 4019 5049 4031 5083
rect 3973 5043 4031 5049
rect 5905 5083 5963 5089
rect 5905 5049 5917 5083
rect 5951 5049 5963 5083
rect 5905 5043 5963 5049
rect 1820 4984 3648 5012
rect 3697 5015 3755 5021
rect 1820 4972 1826 4984
rect 3697 4981 3709 5015
rect 3743 5012 3755 5015
rect 3786 5012 3792 5024
rect 3743 4984 3792 5012
rect 3743 4981 3755 4984
rect 3697 4975 3755 4981
rect 3786 4972 3792 4984
rect 3844 4972 3850 5024
rect 4062 4972 4068 5024
rect 4120 5012 4126 5024
rect 4157 5015 4215 5021
rect 4157 5012 4169 5015
rect 4120 4984 4169 5012
rect 4120 4972 4126 4984
rect 4157 4981 4169 4984
rect 4203 4981 4215 5015
rect 5920 5012 5948 5043
rect 6086 5040 6092 5092
rect 6144 5080 6150 5092
rect 6656 5080 6684 5111
rect 6730 5108 6736 5160
rect 6788 5108 6794 5160
rect 6144 5052 6684 5080
rect 6748 5080 6776 5108
rect 7101 5083 7159 5089
rect 7101 5080 7113 5083
rect 6748 5052 7113 5080
rect 6144 5040 6150 5052
rect 7101 5049 7113 5052
rect 7147 5049 7159 5083
rect 7101 5043 7159 5049
rect 7285 5083 7343 5089
rect 7285 5049 7297 5083
rect 7331 5080 7343 5083
rect 7650 5080 7656 5092
rect 7331 5052 7656 5080
rect 7331 5049 7343 5052
rect 7285 5043 7343 5049
rect 7650 5040 7656 5052
rect 7708 5040 7714 5092
rect 6178 5012 6184 5024
rect 5920 4984 6184 5012
rect 4157 4975 4215 4981
rect 6178 4972 6184 4984
rect 6236 4972 6242 5024
rect 6365 5015 6423 5021
rect 6365 4981 6377 5015
rect 6411 5012 6423 5015
rect 6730 5012 6736 5024
rect 6411 4984 6736 5012
rect 6411 4981 6423 4984
rect 6365 4975 6423 4981
rect 6730 4972 6736 4984
rect 6788 4972 6794 5024
rect 1104 4922 8556 4944
rect 1104 4870 4214 4922
rect 4266 4870 4278 4922
rect 4330 4870 4342 4922
rect 4394 4870 4406 4922
rect 4458 4870 4470 4922
rect 4522 4870 8556 4922
rect 1104 4848 8556 4870
rect 2314 4768 2320 4820
rect 2372 4768 2378 4820
rect 5074 4768 5080 4820
rect 5132 4808 5138 4820
rect 5169 4811 5227 4817
rect 5169 4808 5181 4811
rect 5132 4780 5181 4808
rect 5132 4768 5138 4780
rect 5169 4777 5181 4780
rect 5215 4777 5227 4811
rect 5626 4808 5632 4820
rect 5169 4771 5227 4777
rect 5276 4780 5632 4808
rect 4157 4743 4215 4749
rect 4157 4709 4169 4743
rect 4203 4740 4215 4743
rect 4890 4740 4896 4752
rect 4203 4712 4896 4740
rect 4203 4709 4215 4712
rect 4157 4703 4215 4709
rect 4890 4700 4896 4712
rect 4948 4700 4954 4752
rect 5276 4749 5304 4780
rect 5626 4768 5632 4780
rect 5684 4768 5690 4820
rect 6086 4768 6092 4820
rect 6144 4768 6150 4820
rect 6270 4768 6276 4820
rect 6328 4768 6334 4820
rect 8018 4768 8024 4820
rect 8076 4808 8082 4820
rect 8205 4811 8263 4817
rect 8205 4808 8217 4811
rect 8076 4780 8217 4808
rect 8076 4768 8082 4780
rect 8205 4777 8217 4780
rect 8251 4777 8263 4811
rect 8205 4771 8263 4777
rect 5261 4743 5319 4749
rect 5261 4709 5273 4743
rect 5307 4709 5319 4743
rect 5261 4703 5319 4709
rect 2409 4675 2467 4681
rect 2409 4641 2421 4675
rect 2455 4672 2467 4675
rect 3142 4672 3148 4684
rect 2455 4644 3148 4672
rect 2455 4641 2467 4644
rect 2409 4635 2467 4641
rect 3142 4632 3148 4644
rect 3200 4632 3206 4684
rect 3878 4632 3884 4684
rect 3936 4672 3942 4684
rect 5276 4672 5304 4703
rect 3936 4644 5304 4672
rect 3936 4632 3942 4644
rect 5626 4632 5632 4684
rect 5684 4672 5690 4684
rect 6457 4675 6515 4681
rect 6457 4672 6469 4675
rect 5684 4644 6469 4672
rect 5684 4632 5690 4644
rect 6457 4641 6469 4644
rect 6503 4641 6515 4675
rect 6457 4635 6515 4641
rect 6730 4632 6736 4684
rect 6788 4632 6794 4684
rect 1762 4564 1768 4616
rect 1820 4604 1826 4616
rect 2133 4607 2191 4613
rect 2133 4604 2145 4607
rect 1820 4576 2145 4604
rect 1820 4564 1826 4576
rect 2133 4573 2145 4576
rect 2179 4573 2191 4607
rect 2133 4567 2191 4573
rect 2222 4564 2228 4616
rect 2280 4564 2286 4616
rect 3786 4564 3792 4616
rect 3844 4564 3850 4616
rect 4062 4564 4068 4616
rect 4120 4564 4126 4616
rect 4249 4607 4307 4613
rect 4249 4573 4261 4607
rect 4295 4573 4307 4607
rect 4249 4567 4307 4573
rect 3970 4496 3976 4548
rect 4028 4536 4034 4548
rect 4264 4536 4292 4567
rect 4338 4564 4344 4616
rect 4396 4604 4402 4616
rect 4433 4607 4491 4613
rect 4433 4604 4445 4607
rect 4396 4576 4445 4604
rect 4396 4564 4402 4576
rect 4433 4573 4445 4576
rect 4479 4573 4491 4607
rect 4433 4567 4491 4573
rect 5258 4564 5264 4616
rect 5316 4604 5322 4616
rect 5721 4607 5779 4613
rect 5721 4604 5733 4607
rect 5316 4576 5733 4604
rect 5316 4564 5322 4576
rect 5721 4573 5733 4576
rect 5767 4604 5779 4607
rect 6181 4607 6239 4613
rect 6181 4604 6193 4607
rect 5767 4576 6193 4604
rect 5767 4573 5779 4576
rect 5721 4567 5779 4573
rect 6181 4573 6193 4576
rect 6227 4573 6239 4607
rect 6181 4567 6239 4573
rect 6365 4607 6423 4613
rect 6365 4573 6377 4607
rect 6411 4573 6423 4607
rect 6365 4567 6423 4573
rect 4028 4508 4292 4536
rect 4028 4496 4034 4508
rect 5534 4496 5540 4548
rect 5592 4536 5598 4548
rect 5629 4539 5687 4545
rect 5629 4536 5641 4539
rect 5592 4508 5641 4536
rect 5592 4496 5598 4508
rect 5629 4505 5641 4508
rect 5675 4505 5687 4539
rect 5629 4499 5687 4505
rect 5905 4539 5963 4545
rect 5905 4505 5917 4539
rect 5951 4536 5963 4539
rect 6380 4536 6408 4567
rect 5951 4508 6408 4536
rect 5951 4505 5963 4508
rect 5905 4499 5963 4505
rect 4890 4428 4896 4480
rect 4948 4468 4954 4480
rect 5920 4468 5948 4499
rect 7374 4496 7380 4548
rect 7432 4496 7438 4548
rect 4948 4440 5948 4468
rect 4948 4428 4954 4440
rect 1104 4378 8556 4400
rect 1104 4326 4874 4378
rect 4926 4326 4938 4378
rect 4990 4326 5002 4378
rect 5054 4326 5066 4378
rect 5118 4326 5130 4378
rect 5182 4326 8556 4378
rect 1104 4304 8556 4326
rect 2133 4267 2191 4273
rect 2133 4233 2145 4267
rect 2179 4264 2191 4267
rect 2222 4264 2228 4276
rect 2179 4236 2228 4264
rect 2179 4233 2191 4236
rect 2133 4227 2191 4233
rect 2222 4224 2228 4236
rect 2280 4224 2286 4276
rect 4338 4224 4344 4276
rect 4396 4224 4402 4276
rect 5534 4224 5540 4276
rect 5592 4264 5598 4276
rect 6178 4264 6184 4276
rect 5592 4236 6184 4264
rect 5592 4224 5598 4236
rect 6178 4224 6184 4236
rect 6236 4224 6242 4276
rect 6638 4264 6644 4276
rect 6288 4236 6644 4264
rect 1762 4196 1768 4208
rect 1596 4168 1768 4196
rect 1596 4137 1624 4168
rect 1762 4156 1768 4168
rect 1820 4156 1826 4208
rect 3329 4199 3387 4205
rect 3329 4165 3341 4199
rect 3375 4196 3387 4199
rect 4356 4196 4384 4224
rect 6288 4196 6316 4236
rect 6638 4224 6644 4236
rect 6696 4224 6702 4276
rect 3375 4168 4384 4196
rect 5184 4168 6316 4196
rect 3375 4165 3387 4168
rect 3329 4159 3387 4165
rect 1581 4131 1639 4137
rect 1581 4097 1593 4131
rect 1627 4097 1639 4131
rect 2041 4131 2099 4137
rect 2041 4128 2053 4131
rect 1581 4091 1639 4097
rect 1688 4100 2053 4128
rect 1688 4072 1716 4100
rect 2041 4097 2053 4100
rect 2087 4128 2099 4131
rect 2682 4128 2688 4140
rect 2087 4100 2688 4128
rect 2087 4097 2099 4100
rect 2041 4091 2099 4097
rect 2682 4088 2688 4100
rect 2740 4088 2746 4140
rect 2866 4088 2872 4140
rect 2924 4128 2930 4140
rect 3142 4128 3148 4140
rect 2924 4100 3148 4128
rect 2924 4088 2930 4100
rect 3142 4088 3148 4100
rect 3200 4088 3206 4140
rect 3620 4137 3648 4168
rect 3513 4131 3571 4137
rect 3513 4097 3525 4131
rect 3559 4097 3571 4131
rect 3513 4091 3571 4097
rect 3605 4131 3663 4137
rect 3605 4097 3617 4131
rect 3651 4097 3663 4131
rect 3605 4091 3663 4097
rect 3789 4131 3847 4137
rect 3789 4097 3801 4131
rect 3835 4128 3847 4131
rect 3970 4128 3976 4140
rect 3835 4100 3976 4128
rect 3835 4097 3847 4100
rect 3789 4091 3847 4097
rect 1670 4020 1676 4072
rect 1728 4020 1734 4072
rect 1949 4063 2007 4069
rect 1949 4029 1961 4063
rect 1995 4060 2007 4063
rect 3528 4060 3556 4091
rect 3804 4060 3832 4091
rect 3970 4088 3976 4100
rect 4028 4088 4034 4140
rect 5184 4137 5212 4168
rect 6362 4156 6368 4208
rect 6420 4156 6426 4208
rect 4525 4131 4583 4137
rect 4525 4097 4537 4131
rect 4571 4128 4583 4131
rect 5169 4131 5227 4137
rect 5169 4128 5181 4131
rect 4571 4100 4660 4128
rect 4571 4097 4583 4100
rect 4525 4091 4583 4097
rect 4632 4072 4660 4100
rect 4724 4100 5181 4128
rect 1995 4032 3832 4060
rect 1995 4029 2007 4032
rect 1949 4023 2007 4029
rect 4614 4020 4620 4072
rect 4672 4020 4678 4072
rect 2590 3952 2596 4004
rect 2648 3992 2654 4004
rect 4724 3992 4752 4100
rect 5169 4097 5181 4100
rect 5215 4097 5227 4131
rect 5169 4091 5227 4097
rect 5537 4131 5595 4137
rect 5537 4097 5549 4131
rect 5583 4128 5595 4131
rect 5626 4128 5632 4140
rect 5583 4100 5632 4128
rect 5583 4097 5595 4100
rect 5537 4091 5595 4097
rect 5626 4088 5632 4100
rect 5684 4088 5690 4140
rect 6656 4137 6684 4224
rect 6549 4131 6607 4137
rect 6549 4097 6561 4131
rect 6595 4097 6607 4131
rect 6549 4091 6607 4097
rect 6641 4131 6699 4137
rect 6641 4097 6653 4131
rect 6687 4097 6699 4131
rect 6641 4091 6699 4097
rect 4801 4063 4859 4069
rect 4801 4029 4813 4063
rect 4847 4060 4859 4063
rect 4893 4063 4951 4069
rect 4893 4060 4905 4063
rect 4847 4032 4905 4060
rect 4847 4029 4859 4032
rect 4801 4023 4859 4029
rect 4893 4029 4905 4032
rect 4939 4060 4951 4063
rect 5994 4060 6000 4072
rect 4939 4032 6000 4060
rect 4939 4029 4951 4032
rect 4893 4023 4951 4029
rect 5994 4020 6000 4032
rect 6052 4020 6058 4072
rect 6564 4060 6592 4091
rect 7190 4060 7196 4072
rect 6564 4032 7196 4060
rect 7190 4020 7196 4032
rect 7248 4060 7254 4072
rect 8110 4060 8116 4072
rect 7248 4032 8116 4060
rect 7248 4020 7254 4032
rect 8110 4020 8116 4032
rect 8168 4020 8174 4072
rect 2648 3964 4752 3992
rect 2648 3952 2654 3964
rect 3694 3884 3700 3936
rect 3752 3884 3758 3936
rect 4709 3927 4767 3933
rect 4709 3893 4721 3927
rect 4755 3924 4767 3927
rect 4982 3924 4988 3936
rect 4755 3896 4988 3924
rect 4755 3893 4767 3896
rect 4709 3887 4767 3893
rect 4982 3884 4988 3896
rect 5040 3884 5046 3936
rect 5353 3927 5411 3933
rect 5353 3893 5365 3927
rect 5399 3924 5411 3927
rect 5442 3924 5448 3936
rect 5399 3896 5448 3924
rect 5399 3893 5411 3896
rect 5353 3887 5411 3893
rect 5442 3884 5448 3896
rect 5500 3884 5506 3936
rect 6270 3884 6276 3936
rect 6328 3924 6334 3936
rect 6365 3927 6423 3933
rect 6365 3924 6377 3927
rect 6328 3896 6377 3924
rect 6328 3884 6334 3896
rect 6365 3893 6377 3896
rect 6411 3893 6423 3927
rect 6365 3887 6423 3893
rect 1104 3834 8556 3856
rect 1104 3782 4214 3834
rect 4266 3782 4278 3834
rect 4330 3782 4342 3834
rect 4394 3782 4406 3834
rect 4458 3782 4470 3834
rect 4522 3782 8556 3834
rect 1104 3760 8556 3782
rect 842 3612 848 3664
rect 900 3652 906 3664
rect 1397 3655 1455 3661
rect 1397 3652 1409 3655
rect 900 3624 1409 3652
rect 900 3612 906 3624
rect 1397 3621 1409 3624
rect 1443 3621 1455 3655
rect 1397 3615 1455 3621
rect 4433 3655 4491 3661
rect 4433 3621 4445 3655
rect 4479 3652 4491 3655
rect 4614 3652 4620 3664
rect 4479 3624 4620 3652
rect 4479 3621 4491 3624
rect 4433 3615 4491 3621
rect 4614 3612 4620 3624
rect 4672 3612 4678 3664
rect 2866 3544 2872 3596
rect 2924 3544 2930 3596
rect 2961 3587 3019 3593
rect 2961 3553 2973 3587
rect 3007 3584 3019 3587
rect 3694 3584 3700 3596
rect 3007 3556 3700 3584
rect 3007 3553 3019 3556
rect 2961 3547 3019 3553
rect 3694 3544 3700 3556
rect 3752 3544 3758 3596
rect 4801 3587 4859 3593
rect 4801 3584 4813 3587
rect 4080 3556 4813 3584
rect 1581 3519 1639 3525
rect 1581 3485 1593 3519
rect 1627 3516 1639 3519
rect 1670 3516 1676 3528
rect 1627 3488 1676 3516
rect 1627 3485 1639 3488
rect 1581 3479 1639 3485
rect 1670 3476 1676 3488
rect 1728 3476 1734 3528
rect 2590 3476 2596 3528
rect 2648 3516 2654 3528
rect 3053 3519 3111 3525
rect 3053 3516 3065 3519
rect 2648 3488 3065 3516
rect 2648 3476 2654 3488
rect 3053 3485 3065 3488
rect 3099 3485 3111 3519
rect 3053 3479 3111 3485
rect 3142 3476 3148 3528
rect 3200 3476 3206 3528
rect 3878 3476 3884 3528
rect 3936 3516 3942 3528
rect 4080 3525 4108 3556
rect 4801 3553 4813 3556
rect 4847 3553 4859 3587
rect 4801 3547 4859 3553
rect 4982 3544 4988 3596
rect 5040 3584 5046 3596
rect 5077 3587 5135 3593
rect 5077 3584 5089 3587
rect 5040 3556 5089 3584
rect 5040 3544 5046 3556
rect 5077 3553 5089 3556
rect 5123 3584 5135 3587
rect 5718 3584 5724 3596
rect 5123 3556 5724 3584
rect 5123 3553 5135 3556
rect 5077 3547 5135 3553
rect 5718 3544 5724 3556
rect 5776 3544 5782 3596
rect 4065 3519 4123 3525
rect 4065 3516 4077 3519
rect 3936 3488 4077 3516
rect 3936 3476 3942 3488
rect 4065 3485 4077 3488
rect 4111 3485 4123 3519
rect 4065 3479 4123 3485
rect 4154 3476 4160 3528
rect 4212 3516 4218 3528
rect 4709 3519 4767 3525
rect 4709 3516 4721 3519
rect 4212 3488 4721 3516
rect 4212 3476 4218 3488
rect 4709 3485 4721 3488
rect 4755 3516 4767 3519
rect 5258 3516 5264 3528
rect 4755 3488 5264 3516
rect 4755 3485 4767 3488
rect 4709 3479 4767 3485
rect 5258 3476 5264 3488
rect 5316 3476 5322 3528
rect 5445 3519 5503 3525
rect 5445 3485 5457 3519
rect 5491 3516 5503 3519
rect 5810 3516 5816 3528
rect 5491 3488 5816 3516
rect 5491 3485 5503 3488
rect 5445 3479 5503 3485
rect 5810 3476 5816 3488
rect 5868 3476 5874 3528
rect 7374 3476 7380 3528
rect 7432 3476 7438 3528
rect 7466 3476 7472 3528
rect 7524 3476 7530 3528
rect 2498 3408 2504 3460
rect 2556 3448 2562 3460
rect 4338 3448 4344 3460
rect 2556 3420 4344 3448
rect 2556 3408 2562 3420
rect 4338 3408 4344 3420
rect 4396 3448 4402 3460
rect 7392 3448 7420 3476
rect 4396 3420 7420 3448
rect 4396 3408 4402 3420
rect 2685 3383 2743 3389
rect 2685 3349 2697 3383
rect 2731 3380 2743 3383
rect 2958 3380 2964 3392
rect 2731 3352 2964 3380
rect 2731 3349 2743 3352
rect 2685 3343 2743 3349
rect 2958 3340 2964 3352
rect 3016 3340 3022 3392
rect 6730 3340 6736 3392
rect 6788 3340 6794 3392
rect 7374 3340 7380 3392
rect 7432 3340 7438 3392
rect 1104 3290 8556 3312
rect 1104 3238 4874 3290
rect 4926 3238 4938 3290
rect 4990 3238 5002 3290
rect 5054 3238 5066 3290
rect 5118 3238 5130 3290
rect 5182 3238 8556 3290
rect 1104 3216 8556 3238
rect 1489 3179 1547 3185
rect 1489 3145 1501 3179
rect 1535 3176 1547 3179
rect 1670 3176 1676 3188
rect 1535 3148 1676 3176
rect 1535 3145 1547 3148
rect 1489 3139 1547 3145
rect 1670 3136 1676 3148
rect 1728 3136 1734 3188
rect 3252 3148 5120 3176
rect 2498 3068 2504 3120
rect 2556 3068 2562 3120
rect 2958 3068 2964 3120
rect 3016 3068 3022 3120
rect 3252 3049 3280 3148
rect 4338 3068 4344 3120
rect 4396 3068 4402 3120
rect 5092 3108 5120 3148
rect 8110 3136 8116 3188
rect 8168 3176 8174 3188
rect 8205 3179 8263 3185
rect 8205 3176 8217 3179
rect 8168 3148 8217 3176
rect 8168 3136 8174 3148
rect 8205 3145 8217 3148
rect 8251 3145 8263 3179
rect 8205 3139 8263 3145
rect 5626 3108 5632 3120
rect 5092 3080 5632 3108
rect 5092 3049 5120 3080
rect 5626 3068 5632 3080
rect 5684 3108 5690 3120
rect 6730 3108 6736 3120
rect 5684 3080 6736 3108
rect 5684 3068 5690 3080
rect 3237 3043 3295 3049
rect 3237 3009 3249 3043
rect 3283 3009 3295 3043
rect 3237 3003 3295 3009
rect 5077 3043 5135 3049
rect 5077 3009 5089 3043
rect 5123 3009 5135 3043
rect 5077 3003 5135 3009
rect 5169 3043 5227 3049
rect 5169 3009 5181 3043
rect 5215 3040 5227 3043
rect 5258 3040 5264 3052
rect 5215 3012 5264 3040
rect 5215 3009 5227 3012
rect 5169 3003 5227 3009
rect 5258 3000 5264 3012
rect 5316 3000 5322 3052
rect 5350 3000 5356 3052
rect 5408 3000 5414 3052
rect 5445 3043 5503 3049
rect 5445 3009 5457 3043
rect 5491 3009 5503 3043
rect 5445 3003 5503 3009
rect 3329 2975 3387 2981
rect 3329 2941 3341 2975
rect 3375 2972 3387 2975
rect 4154 2972 4160 2984
rect 3375 2944 4160 2972
rect 3375 2941 3387 2944
rect 3329 2935 3387 2941
rect 4154 2932 4160 2944
rect 4212 2932 4218 2984
rect 4798 2932 4804 2984
rect 4856 2932 4862 2984
rect 4614 2796 4620 2848
rect 4672 2836 4678 2848
rect 5460 2836 5488 3003
rect 5534 3000 5540 3052
rect 5592 3000 5598 3052
rect 5718 3000 5724 3052
rect 5776 3040 5782 3052
rect 5813 3043 5871 3049
rect 5813 3040 5825 3043
rect 5776 3012 5825 3040
rect 5776 3000 5782 3012
rect 5813 3009 5825 3012
rect 5859 3009 5871 3043
rect 5813 3003 5871 3009
rect 5994 3000 6000 3052
rect 6052 3000 6058 3052
rect 6472 3049 6500 3080
rect 6730 3068 6736 3080
rect 6788 3068 6794 3120
rect 7282 3068 7288 3120
rect 7340 3068 7346 3120
rect 6457 3043 6515 3049
rect 6457 3009 6469 3043
rect 6503 3009 6515 3043
rect 6457 3003 6515 3009
rect 6270 2932 6276 2984
rect 6328 2972 6334 2984
rect 6733 2975 6791 2981
rect 6733 2972 6745 2975
rect 6328 2944 6745 2972
rect 6328 2932 6334 2944
rect 6733 2941 6745 2944
rect 6779 2941 6791 2975
rect 6733 2935 6791 2941
rect 5626 2836 5632 2848
rect 4672 2808 5632 2836
rect 4672 2796 4678 2808
rect 5626 2796 5632 2808
rect 5684 2796 5690 2848
rect 5718 2796 5724 2848
rect 5776 2796 5782 2848
rect 5902 2796 5908 2848
rect 5960 2796 5966 2848
rect 1104 2746 8556 2768
rect 1104 2694 4214 2746
rect 4266 2694 4278 2746
rect 4330 2694 4342 2746
rect 4394 2694 4406 2746
rect 4458 2694 4470 2746
rect 4522 2694 8556 2746
rect 1104 2672 8556 2694
rect 3142 2592 3148 2644
rect 3200 2592 3206 2644
rect 3234 2592 3240 2644
rect 3292 2632 3298 2644
rect 4614 2632 4620 2644
rect 3292 2604 4620 2632
rect 3292 2592 3298 2604
rect 4614 2592 4620 2604
rect 4672 2592 4678 2644
rect 4798 2592 4804 2644
rect 4856 2632 4862 2644
rect 4985 2635 5043 2641
rect 4985 2632 4997 2635
rect 4856 2604 4997 2632
rect 4856 2592 4862 2604
rect 4985 2601 4997 2604
rect 5031 2601 5043 2635
rect 4985 2595 5043 2601
rect 5534 2592 5540 2644
rect 5592 2632 5598 2644
rect 5721 2635 5779 2641
rect 5721 2632 5733 2635
rect 5592 2604 5733 2632
rect 5592 2592 5598 2604
rect 5721 2601 5733 2604
rect 5767 2601 5779 2635
rect 5721 2595 5779 2601
rect 6362 2592 6368 2644
rect 6420 2592 6426 2644
rect 6638 2632 6644 2644
rect 6472 2604 6644 2632
rect 3252 2564 3280 2592
rect 2884 2536 3280 2564
rect 1670 2388 1676 2440
rect 1728 2428 1734 2440
rect 2884 2437 2912 2536
rect 5626 2524 5632 2576
rect 5684 2564 5690 2576
rect 6472 2564 6500 2604
rect 6638 2592 6644 2604
rect 6696 2592 6702 2644
rect 7466 2592 7472 2644
rect 7524 2592 7530 2644
rect 7834 2592 7840 2644
rect 7892 2592 7898 2644
rect 5684 2536 6500 2564
rect 5684 2524 5690 2536
rect 6546 2524 6552 2576
rect 6604 2564 6610 2576
rect 7374 2564 7380 2576
rect 6604 2536 7380 2564
rect 6604 2524 6610 2536
rect 7374 2524 7380 2536
rect 7432 2524 7438 2576
rect 3234 2456 3240 2508
rect 3292 2496 3298 2508
rect 5258 2496 5264 2508
rect 3292 2468 3556 2496
rect 3292 2456 3298 2468
rect 3528 2437 3556 2468
rect 4816 2468 5264 2496
rect 4816 2437 4844 2468
rect 5258 2456 5264 2468
rect 5316 2456 5322 2508
rect 5718 2496 5724 2508
rect 5368 2468 5724 2496
rect 2593 2431 2651 2437
rect 2593 2428 2605 2431
rect 1728 2400 2605 2428
rect 1728 2388 1734 2400
rect 2593 2397 2605 2400
rect 2639 2397 2651 2431
rect 2593 2391 2651 2397
rect 2869 2431 2927 2437
rect 2869 2397 2881 2431
rect 2915 2397 2927 2431
rect 2869 2391 2927 2397
rect 2961 2431 3019 2437
rect 2961 2397 2973 2431
rect 3007 2428 3019 2431
rect 3513 2431 3571 2437
rect 3007 2400 3188 2428
rect 3007 2397 3019 2400
rect 2961 2391 3019 2397
rect 2774 2320 2780 2372
rect 2832 2320 2838 2372
rect 3160 2292 3188 2400
rect 3513 2397 3525 2431
rect 3559 2397 3571 2431
rect 3513 2391 3571 2397
rect 4801 2431 4859 2437
rect 4801 2397 4813 2431
rect 4847 2397 4859 2431
rect 4801 2391 4859 2397
rect 5169 2431 5227 2437
rect 5169 2397 5181 2431
rect 5215 2428 5227 2431
rect 5368 2428 5396 2468
rect 5718 2456 5724 2468
rect 5776 2456 5782 2508
rect 5994 2456 6000 2508
rect 6052 2496 6058 2508
rect 7101 2499 7159 2505
rect 7101 2496 7113 2499
rect 6052 2468 7113 2496
rect 6052 2456 6058 2468
rect 5215 2400 5396 2428
rect 5215 2397 5227 2400
rect 5169 2391 5227 2397
rect 5442 2388 5448 2440
rect 5500 2388 5506 2440
rect 5537 2431 5595 2437
rect 5537 2397 5549 2431
rect 5583 2397 5595 2431
rect 5537 2391 5595 2397
rect 5258 2320 5264 2372
rect 5316 2360 5322 2372
rect 5552 2360 5580 2391
rect 6546 2388 6552 2440
rect 6604 2388 6610 2440
rect 6638 2388 6644 2440
rect 6696 2388 6702 2440
rect 6932 2437 6960 2468
rect 7101 2465 7113 2468
rect 7147 2465 7159 2499
rect 7101 2459 7159 2465
rect 7208 2468 7696 2496
rect 7208 2440 7236 2468
rect 6917 2431 6975 2437
rect 6917 2397 6929 2431
rect 6963 2397 6975 2431
rect 6917 2391 6975 2397
rect 7190 2388 7196 2440
rect 7248 2388 7254 2440
rect 7668 2437 7696 2468
rect 7285 2431 7343 2437
rect 7285 2397 7297 2431
rect 7331 2397 7343 2431
rect 7285 2391 7343 2397
rect 7653 2431 7711 2437
rect 7653 2397 7665 2431
rect 7699 2397 7711 2431
rect 7653 2391 7711 2397
rect 5316 2332 5580 2360
rect 5316 2320 5322 2332
rect 5626 2320 5632 2372
rect 5684 2360 5690 2372
rect 6733 2363 6791 2369
rect 6733 2360 6745 2363
rect 5684 2332 6745 2360
rect 5684 2320 5690 2332
rect 6733 2329 6745 2332
rect 6779 2329 6791 2363
rect 7300 2360 7328 2391
rect 8202 2388 8208 2440
rect 8260 2388 8266 2440
rect 6733 2323 6791 2329
rect 6840 2332 7328 2360
rect 3329 2295 3387 2301
rect 3329 2292 3341 2295
rect 3160 2264 3341 2292
rect 3329 2261 3341 2264
rect 3375 2261 3387 2295
rect 3329 2255 3387 2261
rect 4522 2252 4528 2304
rect 4580 2292 4586 2304
rect 4617 2295 4675 2301
rect 4617 2292 4629 2295
rect 4580 2264 4629 2292
rect 4580 2252 4586 2264
rect 4617 2261 4629 2264
rect 4663 2261 4675 2295
rect 4617 2255 4675 2261
rect 5353 2295 5411 2301
rect 5353 2261 5365 2295
rect 5399 2292 5411 2295
rect 5902 2292 5908 2304
rect 5399 2264 5908 2292
rect 5399 2261 5411 2264
rect 5353 2255 5411 2261
rect 5902 2252 5908 2264
rect 5960 2252 5966 2304
rect 6454 2252 6460 2304
rect 6512 2292 6518 2304
rect 6840 2292 6868 2332
rect 6512 2264 6868 2292
rect 6512 2252 6518 2264
rect 7282 2252 7288 2304
rect 7340 2292 7346 2304
rect 8021 2295 8079 2301
rect 8021 2292 8033 2295
rect 7340 2264 8033 2292
rect 7340 2252 7346 2264
rect 8021 2261 8033 2264
rect 8067 2261 8079 2295
rect 8021 2255 8079 2261
rect 1104 2202 8556 2224
rect 1104 2150 4874 2202
rect 4926 2150 4938 2202
rect 4990 2150 5002 2202
rect 5054 2150 5066 2202
rect 5118 2150 5130 2202
rect 5182 2150 8556 2202
rect 1104 2128 8556 2150
rect 2774 2048 2780 2100
rect 2832 2088 2838 2100
rect 5350 2088 5356 2100
rect 2832 2060 5356 2088
rect 2832 2048 2838 2060
rect 5350 2048 5356 2060
rect 5408 2048 5414 2100
<< via1 >>
rect 4214 9222 4266 9274
rect 4278 9222 4330 9274
rect 4342 9222 4394 9274
rect 4406 9222 4458 9274
rect 4470 9222 4522 9274
rect 4620 9163 4672 9172
rect 4620 9129 4629 9163
rect 4629 9129 4663 9163
rect 4663 9129 4672 9163
rect 4620 9120 4672 9129
rect 4804 8959 4856 8968
rect 4804 8925 4813 8959
rect 4813 8925 4847 8959
rect 4847 8925 4856 8959
rect 4804 8916 4856 8925
rect 5172 8916 5224 8968
rect 5264 8823 5316 8832
rect 5264 8789 5273 8823
rect 5273 8789 5307 8823
rect 5307 8789 5316 8823
rect 5264 8780 5316 8789
rect 4874 8678 4926 8730
rect 4938 8678 4990 8730
rect 5002 8678 5054 8730
rect 5066 8678 5118 8730
rect 5130 8678 5182 8730
rect 5632 8619 5684 8628
rect 5632 8585 5641 8619
rect 5641 8585 5675 8619
rect 5675 8585 5684 8619
rect 5632 8576 5684 8585
rect 1584 8483 1636 8492
rect 1584 8449 1593 8483
rect 1593 8449 1627 8483
rect 1627 8449 1636 8483
rect 1584 8440 1636 8449
rect 2044 8483 2096 8492
rect 2044 8449 2053 8483
rect 2053 8449 2087 8483
rect 2087 8449 2096 8483
rect 2044 8440 2096 8449
rect 4528 8508 4580 8560
rect 1400 8347 1452 8356
rect 1400 8313 1409 8347
rect 1409 8313 1443 8347
rect 1443 8313 1452 8347
rect 1400 8304 1452 8313
rect 4344 8483 4396 8492
rect 4344 8449 4353 8483
rect 4353 8449 4387 8483
rect 4387 8449 4396 8483
rect 4344 8440 4396 8449
rect 4528 8372 4580 8424
rect 4988 8415 5040 8424
rect 4988 8381 4997 8415
rect 4997 8381 5031 8415
rect 5031 8381 5040 8415
rect 4988 8372 5040 8381
rect 5908 8304 5960 8356
rect 2780 8279 2832 8288
rect 2780 8245 2789 8279
rect 2789 8245 2823 8279
rect 2823 8245 2832 8279
rect 2780 8236 2832 8245
rect 4344 8236 4396 8288
rect 5448 8236 5500 8288
rect 4214 8134 4266 8186
rect 4278 8134 4330 8186
rect 4342 8134 4394 8186
rect 4406 8134 4458 8186
rect 4470 8134 4522 8186
rect 4344 7939 4396 7948
rect 4344 7905 4353 7939
rect 4353 7905 4387 7939
rect 4387 7905 4396 7939
rect 4344 7896 4396 7905
rect 4436 7939 4488 7948
rect 4436 7905 4445 7939
rect 4445 7905 4479 7939
rect 4479 7905 4488 7939
rect 4436 7896 4488 7905
rect 848 7828 900 7880
rect 2688 7871 2740 7880
rect 2688 7837 2697 7871
rect 2697 7837 2731 7871
rect 2731 7837 2740 7871
rect 2688 7828 2740 7837
rect 2780 7828 2832 7880
rect 5264 7964 5316 8016
rect 4988 7896 5040 7948
rect 5172 7828 5224 7880
rect 5632 7896 5684 7948
rect 6000 7939 6052 7948
rect 6000 7905 6009 7939
rect 6009 7905 6043 7939
rect 6043 7905 6052 7939
rect 6000 7896 6052 7905
rect 2596 7760 2648 7812
rect 4436 7760 4488 7812
rect 4804 7760 4856 7812
rect 5448 7828 5500 7880
rect 5632 7760 5684 7812
rect 2412 7692 2464 7744
rect 2780 7692 2832 7744
rect 3884 7692 3936 7744
rect 4344 7692 4396 7744
rect 5908 7871 5960 7880
rect 5908 7837 5917 7871
rect 5917 7837 5951 7871
rect 5951 7837 5960 7871
rect 5908 7828 5960 7837
rect 6828 7828 6880 7880
rect 6276 7735 6328 7744
rect 6276 7701 6285 7735
rect 6285 7701 6319 7735
rect 6319 7701 6328 7735
rect 6276 7692 6328 7701
rect 8208 7735 8260 7744
rect 8208 7701 8217 7735
rect 8217 7701 8251 7735
rect 8251 7701 8260 7735
rect 8208 7692 8260 7701
rect 4874 7590 4926 7642
rect 4938 7590 4990 7642
rect 5002 7590 5054 7642
rect 5066 7590 5118 7642
rect 5130 7590 5182 7642
rect 3240 7488 3292 7540
rect 4804 7488 4856 7540
rect 7288 7488 7340 7540
rect 2780 7420 2832 7472
rect 5816 7352 5868 7404
rect 7288 7395 7340 7404
rect 7288 7361 7297 7395
rect 7297 7361 7331 7395
rect 7331 7361 7340 7395
rect 7288 7352 7340 7361
rect 7472 7352 7524 7404
rect 3148 7327 3200 7336
rect 3148 7293 3157 7327
rect 3157 7293 3191 7327
rect 3191 7293 3200 7327
rect 3148 7284 3200 7293
rect 6000 7284 6052 7336
rect 6828 7284 6880 7336
rect 8208 7395 8260 7404
rect 8208 7361 8217 7395
rect 8217 7361 8251 7395
rect 8251 7361 8260 7395
rect 8208 7352 8260 7361
rect 5264 7216 5316 7268
rect 7472 7216 7524 7268
rect 1584 7148 1636 7200
rect 4068 7148 4120 7200
rect 7104 7148 7156 7200
rect 4214 7046 4266 7098
rect 4278 7046 4330 7098
rect 4342 7046 4394 7098
rect 4406 7046 4458 7098
rect 4470 7046 4522 7098
rect 1768 6987 1820 6996
rect 1768 6953 1777 6987
rect 1777 6953 1811 6987
rect 1811 6953 1820 6987
rect 1768 6944 1820 6953
rect 2044 6944 2096 6996
rect 2688 6944 2740 6996
rect 3884 6944 3936 6996
rect 5632 6944 5684 6996
rect 6828 6944 6880 6996
rect 5908 6876 5960 6928
rect 4068 6808 4120 6860
rect 6736 6851 6788 6860
rect 6736 6817 6745 6851
rect 6745 6817 6779 6851
rect 6779 6817 6788 6851
rect 6736 6808 6788 6817
rect 940 6740 992 6792
rect 1584 6740 1636 6792
rect 2412 6783 2464 6792
rect 2412 6749 2421 6783
rect 2421 6749 2455 6783
rect 2455 6749 2464 6783
rect 2412 6740 2464 6749
rect 5724 6783 5776 6792
rect 5724 6749 5733 6783
rect 5733 6749 5767 6783
rect 5767 6749 5776 6783
rect 5724 6740 5776 6749
rect 6276 6740 6328 6792
rect 2228 6715 2280 6724
rect 2228 6681 2237 6715
rect 2237 6681 2271 6715
rect 2271 6681 2280 6715
rect 2228 6672 2280 6681
rect 3240 6672 3292 6724
rect 2412 6604 2464 6656
rect 6828 6604 6880 6656
rect 7380 6604 7432 6656
rect 4874 6502 4926 6554
rect 4938 6502 4990 6554
rect 5002 6502 5054 6554
rect 5066 6502 5118 6554
rect 5130 6502 5182 6554
rect 848 6264 900 6316
rect 1860 6307 1912 6316
rect 1860 6273 1869 6307
rect 1869 6273 1903 6307
rect 1903 6273 1912 6307
rect 1860 6264 1912 6273
rect 3148 6400 3200 6452
rect 5356 6400 5408 6452
rect 3240 6332 3292 6384
rect 6276 6400 6328 6452
rect 6736 6400 6788 6452
rect 5908 6332 5960 6384
rect 2780 6239 2832 6248
rect 2780 6205 2789 6239
rect 2789 6205 2823 6239
rect 2823 6205 2832 6239
rect 2780 6196 2832 6205
rect 5172 6239 5224 6248
rect 5172 6205 5181 6239
rect 5181 6205 5215 6239
rect 5215 6205 5224 6239
rect 5172 6196 5224 6205
rect 5264 6239 5316 6248
rect 5264 6205 5273 6239
rect 5273 6205 5307 6239
rect 5307 6205 5316 6239
rect 5264 6196 5316 6205
rect 5632 6196 5684 6248
rect 6000 6307 6052 6316
rect 6000 6273 6009 6307
rect 6009 6273 6043 6307
rect 6043 6273 6052 6307
rect 6000 6264 6052 6273
rect 6184 6307 6236 6316
rect 6184 6273 6193 6307
rect 6193 6273 6227 6307
rect 6227 6273 6236 6307
rect 6184 6264 6236 6273
rect 6828 6307 6880 6316
rect 6828 6273 6837 6307
rect 6837 6273 6871 6307
rect 6871 6273 6880 6307
rect 6828 6264 6880 6273
rect 7104 6307 7156 6316
rect 7104 6273 7113 6307
rect 7113 6273 7147 6307
rect 7147 6273 7156 6307
rect 7104 6264 7156 6273
rect 8024 6307 8076 6316
rect 8024 6273 8033 6307
rect 8033 6273 8067 6307
rect 8067 6273 8076 6307
rect 8024 6264 8076 6273
rect 6736 6196 6788 6248
rect 2504 6128 2556 6180
rect 8208 6171 8260 6180
rect 8208 6137 8217 6171
rect 8217 6137 8251 6171
rect 8251 6137 8260 6171
rect 8208 6128 8260 6137
rect 1676 6103 1728 6112
rect 1676 6069 1685 6103
rect 1685 6069 1719 6103
rect 1719 6069 1728 6103
rect 1676 6060 1728 6069
rect 3792 6060 3844 6112
rect 4214 5958 4266 6010
rect 4278 5958 4330 6010
rect 4342 5958 4394 6010
rect 4406 5958 4458 6010
rect 4470 5958 4522 6010
rect 2780 5856 2832 5908
rect 7472 5788 7524 5840
rect 1860 5720 1912 5772
rect 1768 5652 1820 5704
rect 2044 5695 2096 5704
rect 2044 5661 2053 5695
rect 2053 5661 2087 5695
rect 2087 5661 2096 5695
rect 2044 5652 2096 5661
rect 3792 5720 3844 5772
rect 6184 5720 6236 5772
rect 2504 5695 2556 5704
rect 2504 5661 2518 5695
rect 2518 5661 2552 5695
rect 2552 5661 2556 5695
rect 2504 5652 2556 5661
rect 6920 5695 6972 5704
rect 6920 5661 6929 5695
rect 6929 5661 6963 5695
rect 6963 5661 6972 5695
rect 6920 5652 6972 5661
rect 7196 5652 7248 5704
rect 8024 5720 8076 5772
rect 1952 5559 2004 5568
rect 1952 5525 1961 5559
rect 1961 5525 1995 5559
rect 1995 5525 2004 5559
rect 1952 5516 2004 5525
rect 2228 5516 2280 5568
rect 2412 5627 2464 5636
rect 2412 5593 2421 5627
rect 2421 5593 2455 5627
rect 2455 5593 2464 5627
rect 2412 5584 2464 5593
rect 3240 5584 3292 5636
rect 4620 5584 4672 5636
rect 7656 5695 7708 5704
rect 7656 5661 7665 5695
rect 7665 5661 7699 5695
rect 7699 5661 7708 5695
rect 7656 5652 7708 5661
rect 5080 5516 5132 5568
rect 5448 5516 5500 5568
rect 5816 5559 5868 5568
rect 5816 5525 5825 5559
rect 5825 5525 5859 5559
rect 5859 5525 5868 5559
rect 5816 5516 5868 5525
rect 6828 5516 6880 5568
rect 7472 5516 7524 5568
rect 8208 5695 8260 5704
rect 8208 5661 8217 5695
rect 8217 5661 8251 5695
rect 8251 5661 8260 5695
rect 8208 5652 8260 5661
rect 4874 5414 4926 5466
rect 4938 5414 4990 5466
rect 5002 5414 5054 5466
rect 5066 5414 5118 5466
rect 5130 5414 5182 5466
rect 1952 5312 2004 5364
rect 848 5176 900 5228
rect 2320 5219 2372 5228
rect 2320 5185 2329 5219
rect 2329 5185 2363 5219
rect 2363 5185 2372 5219
rect 2320 5176 2372 5185
rect 4896 5312 4948 5364
rect 5356 5312 5408 5364
rect 5724 5312 5776 5364
rect 6920 5312 6972 5364
rect 2044 5083 2096 5092
rect 2044 5049 2053 5083
rect 2053 5049 2087 5083
rect 2087 5049 2096 5083
rect 2044 5040 2096 5049
rect 2596 5108 2648 5160
rect 2780 5108 2832 5160
rect 3792 5176 3844 5228
rect 7288 5244 7340 5296
rect 5080 5219 5132 5228
rect 5080 5185 5089 5219
rect 5089 5185 5123 5219
rect 5123 5185 5132 5219
rect 5080 5176 5132 5185
rect 5172 5219 5224 5228
rect 5172 5185 5181 5219
rect 5181 5185 5215 5219
rect 5215 5185 5224 5219
rect 5172 5176 5224 5185
rect 5632 5176 5684 5228
rect 6828 5219 6880 5228
rect 6828 5185 6837 5219
rect 6837 5185 6871 5219
rect 6871 5185 6880 5219
rect 6828 5176 6880 5185
rect 6920 5176 6972 5228
rect 8208 5219 8260 5228
rect 8208 5185 8217 5219
rect 8217 5185 8251 5219
rect 8251 5185 8260 5219
rect 8208 5176 8260 5185
rect 6276 5108 6328 5160
rect 2412 5040 2464 5092
rect 1768 4972 1820 5024
rect 3884 5040 3936 5092
rect 3792 4972 3844 5024
rect 4068 4972 4120 5024
rect 6092 5040 6144 5092
rect 6736 5151 6788 5160
rect 6736 5117 6745 5151
rect 6745 5117 6779 5151
rect 6779 5117 6788 5151
rect 6736 5108 6788 5117
rect 7656 5040 7708 5092
rect 6184 4972 6236 5024
rect 6736 4972 6788 5024
rect 4214 4870 4266 4922
rect 4278 4870 4330 4922
rect 4342 4870 4394 4922
rect 4406 4870 4458 4922
rect 4470 4870 4522 4922
rect 2320 4811 2372 4820
rect 2320 4777 2329 4811
rect 2329 4777 2363 4811
rect 2363 4777 2372 4811
rect 2320 4768 2372 4777
rect 5080 4768 5132 4820
rect 4896 4700 4948 4752
rect 5632 4768 5684 4820
rect 6092 4811 6144 4820
rect 6092 4777 6101 4811
rect 6101 4777 6135 4811
rect 6135 4777 6144 4811
rect 6092 4768 6144 4777
rect 6276 4811 6328 4820
rect 6276 4777 6285 4811
rect 6285 4777 6319 4811
rect 6319 4777 6328 4811
rect 6276 4768 6328 4777
rect 8024 4768 8076 4820
rect 3148 4632 3200 4684
rect 3884 4632 3936 4684
rect 5632 4632 5684 4684
rect 6736 4675 6788 4684
rect 6736 4641 6745 4675
rect 6745 4641 6779 4675
rect 6779 4641 6788 4675
rect 6736 4632 6788 4641
rect 1768 4564 1820 4616
rect 2228 4607 2280 4616
rect 2228 4573 2237 4607
rect 2237 4573 2271 4607
rect 2271 4573 2280 4607
rect 2228 4564 2280 4573
rect 3792 4607 3844 4616
rect 3792 4573 3801 4607
rect 3801 4573 3835 4607
rect 3835 4573 3844 4607
rect 3792 4564 3844 4573
rect 4068 4607 4120 4616
rect 4068 4573 4077 4607
rect 4077 4573 4111 4607
rect 4111 4573 4120 4607
rect 4068 4564 4120 4573
rect 3976 4496 4028 4548
rect 4344 4564 4396 4616
rect 5264 4564 5316 4616
rect 5540 4496 5592 4548
rect 4896 4428 4948 4480
rect 7380 4496 7432 4548
rect 4874 4326 4926 4378
rect 4938 4326 4990 4378
rect 5002 4326 5054 4378
rect 5066 4326 5118 4378
rect 5130 4326 5182 4378
rect 2228 4224 2280 4276
rect 4344 4267 4396 4276
rect 4344 4233 4353 4267
rect 4353 4233 4387 4267
rect 4387 4233 4396 4267
rect 4344 4224 4396 4233
rect 5540 4224 5592 4276
rect 6184 4224 6236 4276
rect 1768 4156 1820 4208
rect 6644 4224 6696 4276
rect 2688 4088 2740 4140
rect 2872 4088 2924 4140
rect 3148 4131 3200 4140
rect 3148 4097 3157 4131
rect 3157 4097 3191 4131
rect 3191 4097 3200 4131
rect 3148 4088 3200 4097
rect 1676 4063 1728 4072
rect 1676 4029 1685 4063
rect 1685 4029 1719 4063
rect 1719 4029 1728 4063
rect 1676 4020 1728 4029
rect 3976 4088 4028 4140
rect 6368 4199 6420 4208
rect 6368 4165 6377 4199
rect 6377 4165 6411 4199
rect 6411 4165 6420 4199
rect 6368 4156 6420 4165
rect 4620 4020 4672 4072
rect 2596 3952 2648 4004
rect 5632 4088 5684 4140
rect 6000 4020 6052 4072
rect 7196 4020 7248 4072
rect 8116 4020 8168 4072
rect 3700 3927 3752 3936
rect 3700 3893 3709 3927
rect 3709 3893 3743 3927
rect 3743 3893 3752 3927
rect 3700 3884 3752 3893
rect 4988 3927 5040 3936
rect 4988 3893 4997 3927
rect 4997 3893 5031 3927
rect 5031 3893 5040 3927
rect 4988 3884 5040 3893
rect 5448 3884 5500 3936
rect 6276 3884 6328 3936
rect 4214 3782 4266 3834
rect 4278 3782 4330 3834
rect 4342 3782 4394 3834
rect 4406 3782 4458 3834
rect 4470 3782 4522 3834
rect 848 3612 900 3664
rect 4620 3612 4672 3664
rect 2872 3587 2924 3596
rect 2872 3553 2881 3587
rect 2881 3553 2915 3587
rect 2915 3553 2924 3587
rect 2872 3544 2924 3553
rect 3700 3544 3752 3596
rect 1676 3476 1728 3528
rect 2596 3476 2648 3528
rect 3148 3519 3200 3528
rect 3148 3485 3157 3519
rect 3157 3485 3191 3519
rect 3191 3485 3200 3519
rect 3148 3476 3200 3485
rect 3884 3476 3936 3528
rect 4988 3544 5040 3596
rect 5724 3544 5776 3596
rect 4160 3519 4212 3528
rect 4160 3485 4170 3519
rect 4170 3485 4204 3519
rect 4204 3485 4212 3519
rect 4160 3476 4212 3485
rect 5264 3476 5316 3528
rect 5816 3476 5868 3528
rect 7380 3476 7432 3528
rect 7472 3519 7524 3528
rect 7472 3485 7481 3519
rect 7481 3485 7515 3519
rect 7515 3485 7524 3519
rect 7472 3476 7524 3485
rect 2504 3408 2556 3460
rect 4344 3408 4396 3460
rect 2964 3340 3016 3392
rect 6736 3383 6788 3392
rect 6736 3349 6745 3383
rect 6745 3349 6779 3383
rect 6779 3349 6788 3383
rect 6736 3340 6788 3349
rect 7380 3383 7432 3392
rect 7380 3349 7389 3383
rect 7389 3349 7423 3383
rect 7423 3349 7432 3383
rect 7380 3340 7432 3349
rect 4874 3238 4926 3290
rect 4938 3238 4990 3290
rect 5002 3238 5054 3290
rect 5066 3238 5118 3290
rect 5130 3238 5182 3290
rect 1676 3136 1728 3188
rect 2504 3068 2556 3120
rect 2964 3111 3016 3120
rect 2964 3077 2973 3111
rect 2973 3077 3007 3111
rect 3007 3077 3016 3111
rect 2964 3068 3016 3077
rect 4344 3068 4396 3120
rect 8116 3136 8168 3188
rect 5632 3068 5684 3120
rect 5264 3000 5316 3052
rect 5356 3043 5408 3052
rect 5356 3009 5365 3043
rect 5365 3009 5399 3043
rect 5399 3009 5408 3043
rect 5356 3000 5408 3009
rect 4160 2932 4212 2984
rect 4804 2975 4856 2984
rect 4804 2941 4813 2975
rect 4813 2941 4847 2975
rect 4847 2941 4856 2975
rect 4804 2932 4856 2941
rect 4620 2796 4672 2848
rect 5540 3043 5592 3052
rect 5540 3009 5549 3043
rect 5549 3009 5583 3043
rect 5583 3009 5592 3043
rect 5540 3000 5592 3009
rect 5724 3000 5776 3052
rect 6000 3043 6052 3052
rect 6000 3009 6009 3043
rect 6009 3009 6043 3043
rect 6043 3009 6052 3043
rect 6000 3000 6052 3009
rect 6736 3068 6788 3120
rect 7288 3068 7340 3120
rect 6276 2932 6328 2984
rect 5632 2796 5684 2848
rect 5724 2839 5776 2848
rect 5724 2805 5733 2839
rect 5733 2805 5767 2839
rect 5767 2805 5776 2839
rect 5724 2796 5776 2805
rect 5908 2839 5960 2848
rect 5908 2805 5917 2839
rect 5917 2805 5951 2839
rect 5951 2805 5960 2839
rect 5908 2796 5960 2805
rect 4214 2694 4266 2746
rect 4278 2694 4330 2746
rect 4342 2694 4394 2746
rect 4406 2694 4458 2746
rect 4470 2694 4522 2746
rect 3148 2635 3200 2644
rect 3148 2601 3157 2635
rect 3157 2601 3191 2635
rect 3191 2601 3200 2635
rect 3148 2592 3200 2601
rect 3240 2592 3292 2644
rect 4620 2592 4672 2644
rect 4804 2592 4856 2644
rect 5540 2592 5592 2644
rect 6368 2635 6420 2644
rect 6368 2601 6377 2635
rect 6377 2601 6411 2635
rect 6411 2601 6420 2635
rect 6368 2592 6420 2601
rect 1676 2388 1728 2440
rect 5632 2524 5684 2576
rect 6644 2592 6696 2644
rect 7472 2635 7524 2644
rect 7472 2601 7481 2635
rect 7481 2601 7515 2635
rect 7515 2601 7524 2635
rect 7472 2592 7524 2601
rect 7840 2635 7892 2644
rect 7840 2601 7849 2635
rect 7849 2601 7883 2635
rect 7883 2601 7892 2635
rect 7840 2592 7892 2601
rect 6552 2524 6604 2576
rect 7380 2524 7432 2576
rect 3240 2456 3292 2508
rect 5264 2456 5316 2508
rect 2780 2363 2832 2372
rect 2780 2329 2789 2363
rect 2789 2329 2823 2363
rect 2823 2329 2832 2363
rect 2780 2320 2832 2329
rect 5724 2456 5776 2508
rect 6000 2456 6052 2508
rect 5448 2431 5500 2440
rect 5448 2397 5457 2431
rect 5457 2397 5491 2431
rect 5491 2397 5500 2431
rect 5448 2388 5500 2397
rect 5264 2320 5316 2372
rect 6552 2431 6604 2440
rect 6552 2397 6561 2431
rect 6561 2397 6595 2431
rect 6595 2397 6604 2431
rect 6552 2388 6604 2397
rect 6644 2431 6696 2440
rect 6644 2397 6653 2431
rect 6653 2397 6687 2431
rect 6687 2397 6696 2431
rect 6644 2388 6696 2397
rect 7196 2431 7248 2440
rect 7196 2397 7205 2431
rect 7205 2397 7239 2431
rect 7239 2397 7248 2431
rect 7196 2388 7248 2397
rect 5632 2320 5684 2372
rect 8208 2431 8260 2440
rect 8208 2397 8217 2431
rect 8217 2397 8251 2431
rect 8251 2397 8260 2431
rect 8208 2388 8260 2397
rect 4528 2252 4580 2304
rect 5908 2252 5960 2304
rect 6460 2252 6512 2304
rect 7288 2252 7340 2304
rect 4874 2150 4926 2202
rect 4938 2150 4990 2202
rect 5002 2150 5054 2202
rect 5066 2150 5118 2202
rect 5130 2150 5182 2202
rect 2780 2048 2832 2100
rect 5356 2048 5408 2100
<< metal2 >>
rect 4526 11019 4582 11819
rect 5170 11019 5226 11819
rect 4540 10010 4568 11019
rect 4540 9982 4660 10010
rect 4214 9276 4522 9285
rect 4214 9274 4220 9276
rect 4276 9274 4300 9276
rect 4356 9274 4380 9276
rect 4436 9274 4460 9276
rect 4516 9274 4522 9276
rect 4276 9222 4278 9274
rect 4458 9222 4460 9274
rect 4214 9220 4220 9222
rect 4276 9220 4300 9222
rect 4356 9220 4380 9222
rect 4436 9220 4460 9222
rect 4516 9220 4522 9222
rect 4214 9211 4522 9220
rect 4632 9178 4660 9982
rect 4620 9172 4672 9178
rect 4620 9114 4672 9120
rect 5184 8974 5212 11019
rect 4804 8968 4856 8974
rect 4804 8910 4856 8916
rect 5172 8968 5224 8974
rect 5172 8910 5224 8916
rect 4528 8560 4580 8566
rect 4528 8502 4580 8508
rect 4816 8514 4844 8910
rect 5264 8832 5316 8838
rect 5264 8774 5316 8780
rect 4874 8732 5182 8741
rect 4874 8730 4880 8732
rect 4936 8730 4960 8732
rect 5016 8730 5040 8732
rect 5096 8730 5120 8732
rect 5176 8730 5182 8732
rect 4936 8678 4938 8730
rect 5118 8678 5120 8730
rect 4874 8676 4880 8678
rect 4936 8676 4960 8678
rect 5016 8676 5040 8678
rect 5096 8676 5120 8678
rect 5176 8676 5182 8678
rect 4874 8667 5182 8676
rect 1584 8492 1636 8498
rect 1584 8434 1636 8440
rect 2044 8492 2096 8498
rect 2044 8434 2096 8440
rect 4344 8492 4396 8498
rect 4344 8434 4396 8440
rect 1400 8356 1452 8362
rect 1400 8298 1452 8304
rect 1412 8265 1440 8298
rect 1398 8256 1454 8265
rect 1398 8191 1454 8200
rect 848 7880 900 7886
rect 848 7822 900 7828
rect 860 7721 888 7822
rect 846 7712 902 7721
rect 846 7647 902 7656
rect 1596 7206 1624 8434
rect 1584 7200 1636 7206
rect 1584 7142 1636 7148
rect 938 6896 994 6905
rect 938 6831 994 6840
rect 952 6798 980 6831
rect 1596 6798 1624 7142
rect 2056 7002 2084 8434
rect 4356 8294 4384 8434
rect 4540 8430 4568 8502
rect 4816 8486 5028 8514
rect 5000 8430 5028 8486
rect 4528 8424 4580 8430
rect 4528 8366 4580 8372
rect 4988 8424 5040 8430
rect 4988 8366 5040 8372
rect 2780 8288 2832 8294
rect 2780 8230 2832 8236
rect 4344 8288 4396 8294
rect 4344 8230 4396 8236
rect 2792 7886 2820 8230
rect 4214 8188 4522 8197
rect 4214 8186 4220 8188
rect 4276 8186 4300 8188
rect 4356 8186 4380 8188
rect 4436 8186 4460 8188
rect 4516 8186 4522 8188
rect 4276 8134 4278 8186
rect 4458 8134 4460 8186
rect 4214 8132 4220 8134
rect 4276 8132 4300 8134
rect 4356 8132 4380 8134
rect 4436 8132 4460 8134
rect 4516 8132 4522 8134
rect 4214 8123 4522 8132
rect 5000 7954 5028 8366
rect 5276 8022 5304 8774
rect 5632 8628 5684 8634
rect 5632 8570 5684 8576
rect 5448 8288 5500 8294
rect 5448 8230 5500 8236
rect 5264 8016 5316 8022
rect 5264 7958 5316 7964
rect 4344 7948 4396 7954
rect 4344 7890 4396 7896
rect 4436 7948 4488 7954
rect 4436 7890 4488 7896
rect 4988 7948 5040 7954
rect 4988 7890 5040 7896
rect 2688 7880 2740 7886
rect 2688 7822 2740 7828
rect 2780 7880 2832 7886
rect 2780 7822 2832 7828
rect 2596 7812 2648 7818
rect 2596 7754 2648 7760
rect 2412 7744 2464 7750
rect 2412 7686 2464 7692
rect 1768 6996 1820 7002
rect 1768 6938 1820 6944
rect 2044 6996 2096 7002
rect 2044 6938 2096 6944
rect 940 6792 992 6798
rect 940 6734 992 6740
rect 1584 6792 1636 6798
rect 1584 6734 1636 6740
rect 848 6316 900 6322
rect 848 6258 900 6264
rect 860 6089 888 6258
rect 1676 6112 1728 6118
rect 846 6080 902 6089
rect 1676 6054 1728 6060
rect 846 6015 902 6024
rect 1688 5545 1716 6054
rect 1780 5710 1808 6938
rect 2424 6798 2452 7686
rect 2412 6792 2464 6798
rect 2412 6734 2464 6740
rect 2228 6724 2280 6730
rect 2228 6666 2280 6672
rect 1860 6316 1912 6322
rect 1860 6258 1912 6264
rect 1872 5778 1900 6258
rect 1860 5772 1912 5778
rect 1860 5714 1912 5720
rect 1768 5704 1820 5710
rect 1768 5646 1820 5652
rect 2044 5704 2096 5710
rect 2044 5646 2096 5652
rect 1674 5536 1730 5545
rect 1674 5471 1730 5480
rect 848 5228 900 5234
rect 848 5170 900 5176
rect 860 5001 888 5170
rect 1780 5030 1808 5646
rect 1952 5568 2004 5574
rect 1952 5510 2004 5516
rect 1964 5370 1992 5510
rect 1952 5364 2004 5370
rect 1952 5306 2004 5312
rect 2056 5098 2084 5646
rect 2240 5574 2268 6666
rect 2412 6656 2464 6662
rect 2412 6598 2464 6604
rect 2424 5642 2452 6598
rect 2504 6180 2556 6186
rect 2504 6122 2556 6128
rect 2516 5710 2544 6122
rect 2504 5704 2556 5710
rect 2504 5646 2556 5652
rect 2412 5636 2464 5642
rect 2412 5578 2464 5584
rect 2228 5568 2280 5574
rect 2228 5510 2280 5516
rect 2320 5228 2372 5234
rect 2320 5170 2372 5176
rect 2044 5092 2096 5098
rect 2044 5034 2096 5040
rect 1768 5024 1820 5030
rect 846 4992 902 5001
rect 1768 4966 1820 4972
rect 846 4927 902 4936
rect 1780 4622 1808 4966
rect 2332 4826 2360 5170
rect 2424 5098 2452 5578
rect 2608 5166 2636 7754
rect 2700 7002 2728 7822
rect 4356 7750 4384 7890
rect 4448 7818 4476 7890
rect 5460 7886 5488 8230
rect 5644 7954 5672 8570
rect 5908 8356 5960 8362
rect 5908 8298 5960 8304
rect 5632 7948 5684 7954
rect 5632 7890 5684 7896
rect 5920 7886 5948 8298
rect 6000 7948 6052 7954
rect 6000 7890 6052 7896
rect 5172 7880 5224 7886
rect 5448 7880 5500 7886
rect 5224 7840 5304 7868
rect 5172 7822 5224 7828
rect 4436 7812 4488 7818
rect 4436 7754 4488 7760
rect 4804 7812 4856 7818
rect 4804 7754 4856 7760
rect 2780 7744 2832 7750
rect 2780 7686 2832 7692
rect 3884 7744 3936 7750
rect 3884 7686 3936 7692
rect 4344 7744 4396 7750
rect 4344 7686 4396 7692
rect 2792 7478 2820 7686
rect 3240 7540 3292 7546
rect 3240 7482 3292 7488
rect 2780 7472 2832 7478
rect 2780 7414 2832 7420
rect 3148 7336 3200 7342
rect 3148 7278 3200 7284
rect 2688 6996 2740 7002
rect 2688 6938 2740 6944
rect 3160 6458 3188 7278
rect 3252 6730 3280 7482
rect 3896 7002 3924 7686
rect 4816 7546 4844 7754
rect 4874 7644 5182 7653
rect 4874 7642 4880 7644
rect 4936 7642 4960 7644
rect 5016 7642 5040 7644
rect 5096 7642 5120 7644
rect 5176 7642 5182 7644
rect 4936 7590 4938 7642
rect 5118 7590 5120 7642
rect 4874 7588 4880 7590
rect 4936 7588 4960 7590
rect 5016 7588 5040 7590
rect 5096 7588 5120 7590
rect 5176 7588 5182 7590
rect 4874 7579 5182 7588
rect 4804 7540 4856 7546
rect 4804 7482 4856 7488
rect 5276 7274 5304 7840
rect 5368 7840 5448 7868
rect 5264 7268 5316 7274
rect 5264 7210 5316 7216
rect 4068 7200 4120 7206
rect 4068 7142 4120 7148
rect 3884 6996 3936 7002
rect 3884 6938 3936 6944
rect 4080 6866 4108 7142
rect 4214 7100 4522 7109
rect 4214 7098 4220 7100
rect 4276 7098 4300 7100
rect 4356 7098 4380 7100
rect 4436 7098 4460 7100
rect 4516 7098 4522 7100
rect 4276 7046 4278 7098
rect 4458 7046 4460 7098
rect 4214 7044 4220 7046
rect 4276 7044 4300 7046
rect 4356 7044 4380 7046
rect 4436 7044 4460 7046
rect 4516 7044 4522 7046
rect 4214 7035 4522 7044
rect 4068 6860 4120 6866
rect 4068 6802 4120 6808
rect 3240 6724 3292 6730
rect 3240 6666 3292 6672
rect 3148 6452 3200 6458
rect 3148 6394 3200 6400
rect 3252 6390 3280 6666
rect 4874 6556 5182 6565
rect 4874 6554 4880 6556
rect 4936 6554 4960 6556
rect 5016 6554 5040 6556
rect 5096 6554 5120 6556
rect 5176 6554 5182 6556
rect 4936 6502 4938 6554
rect 5118 6502 5120 6554
rect 4874 6500 4880 6502
rect 4936 6500 4960 6502
rect 5016 6500 5040 6502
rect 5096 6500 5120 6502
rect 5176 6500 5182 6502
rect 4874 6491 5182 6500
rect 3240 6384 3292 6390
rect 5276 6338 5304 7210
rect 5368 6458 5396 7840
rect 5448 7822 5500 7828
rect 5908 7880 5960 7886
rect 5908 7822 5960 7828
rect 5632 7812 5684 7818
rect 5632 7754 5684 7760
rect 5644 7002 5672 7754
rect 5816 7404 5868 7410
rect 5816 7346 5868 7352
rect 5632 6996 5684 7002
rect 5632 6938 5684 6944
rect 5724 6792 5776 6798
rect 5724 6734 5776 6740
rect 5356 6452 5408 6458
rect 5356 6394 5408 6400
rect 3240 6326 3292 6332
rect 5092 6310 5304 6338
rect 2780 6248 2832 6254
rect 2780 6190 2832 6196
rect 2792 5914 2820 6190
rect 3792 6112 3844 6118
rect 3792 6054 3844 6060
rect 2780 5908 2832 5914
rect 2780 5850 2832 5856
rect 3804 5778 3832 6054
rect 4214 6012 4522 6021
rect 4214 6010 4220 6012
rect 4276 6010 4300 6012
rect 4356 6010 4380 6012
rect 4436 6010 4460 6012
rect 4516 6010 4522 6012
rect 4276 5958 4278 6010
rect 4458 5958 4460 6010
rect 4214 5956 4220 5958
rect 4276 5956 4300 5958
rect 4356 5956 4380 5958
rect 4436 5956 4460 5958
rect 4516 5956 4522 5958
rect 4214 5947 4522 5956
rect 3792 5772 3844 5778
rect 3792 5714 3844 5720
rect 3240 5636 3292 5642
rect 3240 5578 3292 5584
rect 2596 5160 2648 5166
rect 2780 5160 2832 5166
rect 2596 5102 2648 5108
rect 2700 5108 2780 5114
rect 2700 5102 2832 5108
rect 2412 5092 2464 5098
rect 2412 5034 2464 5040
rect 2320 4820 2372 4826
rect 2320 4762 2372 4768
rect 1768 4616 1820 4622
rect 1768 4558 1820 4564
rect 2228 4616 2280 4622
rect 2228 4558 2280 4564
rect 1780 4214 1808 4558
rect 2240 4282 2268 4558
rect 2228 4276 2280 4282
rect 2228 4218 2280 4224
rect 1768 4208 1820 4214
rect 1768 4150 1820 4156
rect 1676 4072 1728 4078
rect 1676 4014 1728 4020
rect 848 3664 900 3670
rect 846 3632 848 3641
rect 900 3632 902 3641
rect 846 3567 902 3576
rect 1688 3534 1716 4014
rect 2608 4010 2636 5102
rect 2700 5086 2820 5102
rect 2700 4146 2728 5086
rect 3148 4684 3200 4690
rect 3148 4626 3200 4632
rect 3160 4146 3188 4626
rect 2688 4140 2740 4146
rect 2688 4082 2740 4088
rect 2872 4140 2924 4146
rect 2872 4082 2924 4088
rect 3148 4140 3200 4146
rect 3148 4082 3200 4088
rect 2596 4004 2648 4010
rect 2596 3946 2648 3952
rect 2608 3534 2636 3946
rect 2884 3602 2912 4082
rect 2872 3596 2924 3602
rect 2872 3538 2924 3544
rect 1676 3528 1728 3534
rect 1676 3470 1728 3476
rect 2596 3528 2648 3534
rect 2596 3470 2648 3476
rect 3148 3528 3200 3534
rect 3148 3470 3200 3476
rect 1688 3194 1716 3470
rect 2504 3460 2556 3466
rect 2504 3402 2556 3408
rect 1676 3188 1728 3194
rect 1676 3130 1728 3136
rect 1688 2446 1716 3130
rect 2516 3126 2544 3402
rect 2964 3392 3016 3398
rect 2964 3334 3016 3340
rect 2976 3126 3004 3334
rect 2504 3120 2556 3126
rect 2504 3062 2556 3068
rect 2964 3120 3016 3126
rect 2964 3062 3016 3068
rect 3160 2650 3188 3470
rect 3252 2650 3280 5578
rect 3804 5234 3832 5714
rect 4620 5636 4672 5642
rect 4620 5578 4672 5584
rect 3792 5228 3844 5234
rect 3792 5170 3844 5176
rect 3884 5092 3936 5098
rect 3884 5034 3936 5040
rect 3792 5024 3844 5030
rect 3792 4966 3844 4972
rect 3804 4622 3832 4966
rect 3896 4690 3924 5034
rect 4068 5024 4120 5030
rect 4068 4966 4120 4972
rect 3884 4684 3936 4690
rect 3884 4626 3936 4632
rect 3792 4616 3844 4622
rect 3792 4558 3844 4564
rect 3700 3936 3752 3942
rect 3700 3878 3752 3884
rect 3712 3602 3740 3878
rect 3700 3596 3752 3602
rect 3700 3538 3752 3544
rect 3896 3534 3924 4626
rect 4080 4622 4108 4966
rect 4214 4924 4522 4933
rect 4214 4922 4220 4924
rect 4276 4922 4300 4924
rect 4356 4922 4380 4924
rect 4436 4922 4460 4924
rect 4516 4922 4522 4924
rect 4276 4870 4278 4922
rect 4458 4870 4460 4922
rect 4214 4868 4220 4870
rect 4276 4868 4300 4870
rect 4356 4868 4380 4870
rect 4436 4868 4460 4870
rect 4516 4868 4522 4870
rect 4214 4859 4522 4868
rect 4068 4616 4120 4622
rect 4068 4558 4120 4564
rect 4344 4616 4396 4622
rect 4344 4558 4396 4564
rect 3976 4548 4028 4554
rect 3976 4490 4028 4496
rect 3988 4146 4016 4490
rect 4356 4282 4384 4558
rect 4344 4276 4396 4282
rect 4344 4218 4396 4224
rect 4632 4185 4660 5578
rect 5092 5574 5120 6310
rect 5172 6248 5224 6254
rect 5172 6190 5224 6196
rect 5264 6248 5316 6254
rect 5264 6190 5316 6196
rect 5632 6248 5684 6254
rect 5632 6190 5684 6196
rect 5184 5624 5212 6190
rect 5276 5692 5304 6190
rect 5276 5664 5396 5692
rect 5184 5596 5304 5624
rect 5080 5568 5132 5574
rect 5080 5510 5132 5516
rect 4874 5468 5182 5477
rect 4874 5466 4880 5468
rect 4936 5466 4960 5468
rect 5016 5466 5040 5468
rect 5096 5466 5120 5468
rect 5176 5466 5182 5468
rect 4936 5414 4938 5466
rect 5118 5414 5120 5466
rect 4874 5412 4880 5414
rect 4936 5412 4960 5414
rect 5016 5412 5040 5414
rect 5096 5412 5120 5414
rect 5176 5412 5182 5414
rect 4874 5403 5182 5412
rect 4896 5364 4948 5370
rect 4896 5306 4948 5312
rect 4908 4758 4936 5306
rect 5080 5228 5132 5234
rect 5080 5170 5132 5176
rect 5172 5228 5224 5234
rect 5276 5216 5304 5596
rect 5368 5370 5396 5664
rect 5448 5568 5500 5574
rect 5448 5510 5500 5516
rect 5356 5364 5408 5370
rect 5356 5306 5408 5312
rect 5460 5250 5488 5510
rect 5224 5188 5304 5216
rect 5172 5170 5224 5176
rect 5092 4826 5120 5170
rect 5080 4820 5132 4826
rect 5080 4762 5132 4768
rect 4896 4752 4948 4758
rect 4896 4694 4948 4700
rect 4908 4486 4936 4694
rect 5276 4622 5304 5188
rect 5368 5222 5488 5250
rect 5644 5234 5672 6190
rect 5736 5370 5764 6734
rect 5828 5574 5856 7346
rect 6012 7342 6040 7890
rect 6828 7880 6880 7886
rect 6828 7822 6880 7828
rect 6276 7744 6328 7750
rect 6276 7686 6328 7692
rect 6000 7336 6052 7342
rect 6000 7278 6052 7284
rect 5908 6928 5960 6934
rect 5908 6870 5960 6876
rect 5920 6390 5948 6870
rect 5908 6384 5960 6390
rect 5908 6326 5960 6332
rect 6012 6322 6040 7278
rect 6288 6798 6316 7686
rect 6840 7342 6868 7822
rect 8208 7744 8260 7750
rect 8208 7686 8260 7692
rect 8220 7585 8248 7686
rect 8206 7576 8262 7585
rect 7288 7540 7340 7546
rect 8206 7511 8262 7520
rect 7288 7482 7340 7488
rect 7300 7410 7328 7482
rect 7288 7404 7340 7410
rect 7288 7346 7340 7352
rect 7472 7404 7524 7410
rect 7472 7346 7524 7352
rect 8208 7404 8260 7410
rect 8208 7346 8260 7352
rect 6828 7336 6880 7342
rect 6828 7278 6880 7284
rect 6840 7002 6868 7278
rect 7104 7200 7156 7206
rect 7104 7142 7156 7148
rect 6828 6996 6880 7002
rect 6828 6938 6880 6944
rect 6736 6860 6788 6866
rect 6736 6802 6788 6808
rect 6276 6792 6328 6798
rect 6276 6734 6328 6740
rect 6288 6458 6316 6734
rect 6748 6458 6776 6802
rect 6828 6656 6880 6662
rect 6828 6598 6880 6604
rect 6276 6452 6328 6458
rect 6276 6394 6328 6400
rect 6736 6452 6788 6458
rect 6736 6394 6788 6400
rect 6840 6322 6868 6598
rect 7116 6322 7144 7142
rect 6000 6316 6052 6322
rect 6000 6258 6052 6264
rect 6184 6316 6236 6322
rect 6184 6258 6236 6264
rect 6828 6316 6880 6322
rect 6828 6258 6880 6264
rect 7104 6316 7156 6322
rect 7104 6258 7156 6264
rect 6196 5778 6224 6258
rect 6736 6248 6788 6254
rect 6736 6190 6788 6196
rect 6184 5772 6236 5778
rect 6184 5714 6236 5720
rect 5816 5568 5868 5574
rect 5816 5510 5868 5516
rect 5724 5364 5776 5370
rect 5724 5306 5776 5312
rect 5632 5228 5684 5234
rect 5264 4616 5316 4622
rect 5264 4558 5316 4564
rect 4896 4480 4948 4486
rect 4896 4422 4948 4428
rect 4874 4380 5182 4389
rect 4874 4378 4880 4380
rect 4936 4378 4960 4380
rect 5016 4378 5040 4380
rect 5096 4378 5120 4380
rect 5176 4378 5182 4380
rect 4936 4326 4938 4378
rect 5118 4326 5120 4378
rect 4874 4324 4880 4326
rect 4936 4324 4960 4326
rect 5016 4324 5040 4326
rect 5096 4324 5120 4326
rect 5176 4324 5182 4326
rect 4874 4315 5182 4324
rect 4618 4176 4674 4185
rect 3976 4140 4028 4146
rect 4618 4111 4674 4120
rect 3976 4082 4028 4088
rect 4620 4072 4672 4078
rect 4620 4014 4672 4020
rect 4214 3836 4522 3845
rect 4214 3834 4220 3836
rect 4276 3834 4300 3836
rect 4356 3834 4380 3836
rect 4436 3834 4460 3836
rect 4516 3834 4522 3836
rect 4276 3782 4278 3834
rect 4458 3782 4460 3834
rect 4214 3780 4220 3782
rect 4276 3780 4300 3782
rect 4356 3780 4380 3782
rect 4436 3780 4460 3782
rect 4516 3780 4522 3782
rect 4214 3771 4522 3780
rect 4632 3670 4660 4014
rect 4988 3936 5040 3942
rect 4988 3878 5040 3884
rect 4620 3664 4672 3670
rect 4620 3606 4672 3612
rect 5000 3602 5028 3878
rect 4988 3596 5040 3602
rect 4988 3538 5040 3544
rect 3884 3528 3936 3534
rect 3884 3470 3936 3476
rect 4160 3528 4212 3534
rect 4160 3470 4212 3476
rect 5264 3528 5316 3534
rect 5264 3470 5316 3476
rect 4172 2990 4200 3470
rect 4344 3460 4396 3466
rect 4344 3402 4396 3408
rect 4356 3126 4384 3402
rect 4874 3292 5182 3301
rect 4874 3290 4880 3292
rect 4936 3290 4960 3292
rect 5016 3290 5040 3292
rect 5096 3290 5120 3292
rect 5176 3290 5182 3292
rect 4936 3238 4938 3290
rect 5118 3238 5120 3290
rect 4874 3236 4880 3238
rect 4936 3236 4960 3238
rect 5016 3236 5040 3238
rect 5096 3236 5120 3238
rect 5176 3236 5182 3238
rect 4874 3227 5182 3236
rect 4344 3120 4396 3126
rect 4344 3062 4396 3068
rect 5276 3058 5304 3470
rect 5368 3058 5396 5222
rect 5632 5170 5684 5176
rect 5644 4826 5672 5170
rect 5632 4820 5684 4826
rect 5632 4762 5684 4768
rect 5632 4684 5684 4690
rect 5632 4626 5684 4632
rect 5540 4548 5592 4554
rect 5540 4490 5592 4496
rect 5552 4282 5580 4490
rect 5540 4276 5592 4282
rect 5540 4218 5592 4224
rect 5644 4146 5672 4626
rect 5632 4140 5684 4146
rect 5632 4082 5684 4088
rect 5448 3936 5500 3942
rect 5448 3878 5500 3884
rect 5264 3052 5316 3058
rect 5264 2994 5316 3000
rect 5356 3052 5408 3058
rect 5356 2994 5408 3000
rect 4160 2984 4212 2990
rect 4160 2926 4212 2932
rect 4804 2984 4856 2990
rect 4804 2926 4856 2932
rect 4620 2848 4672 2854
rect 4620 2790 4672 2796
rect 4214 2748 4522 2757
rect 4214 2746 4220 2748
rect 4276 2746 4300 2748
rect 4356 2746 4380 2748
rect 4436 2746 4460 2748
rect 4516 2746 4522 2748
rect 4276 2694 4278 2746
rect 4458 2694 4460 2746
rect 4214 2692 4220 2694
rect 4276 2692 4300 2694
rect 4356 2692 4380 2694
rect 4436 2692 4460 2694
rect 4516 2692 4522 2694
rect 4214 2683 4522 2692
rect 4632 2650 4660 2790
rect 4816 2650 4844 2926
rect 3148 2644 3200 2650
rect 3148 2586 3200 2592
rect 3240 2644 3292 2650
rect 3240 2586 3292 2592
rect 4620 2644 4672 2650
rect 4620 2586 4672 2592
rect 4804 2644 4856 2650
rect 4804 2586 4856 2592
rect 5276 2514 5304 2994
rect 3240 2508 3292 2514
rect 3240 2450 3292 2456
rect 5264 2508 5316 2514
rect 5264 2450 5316 2456
rect 1676 2440 1728 2446
rect 1676 2382 1728 2388
rect 2780 2372 2832 2378
rect 2780 2314 2832 2320
rect 2792 2106 2820 2314
rect 2780 2100 2832 2106
rect 2780 2042 2832 2048
rect 3252 800 3280 2450
rect 5264 2372 5316 2378
rect 5264 2314 5316 2320
rect 4528 2304 4580 2310
rect 4528 2246 4580 2252
rect 4540 800 4568 2246
rect 4874 2204 5182 2213
rect 4874 2202 4880 2204
rect 4936 2202 4960 2204
rect 5016 2202 5040 2204
rect 5096 2202 5120 2204
rect 5176 2202 5182 2204
rect 4936 2150 4938 2202
rect 5118 2150 5120 2202
rect 4874 2148 4880 2150
rect 4936 2148 4960 2150
rect 5016 2148 5040 2150
rect 5096 2148 5120 2150
rect 5176 2148 5182 2150
rect 4874 2139 5182 2148
rect 5276 1306 5304 2314
rect 5368 2258 5396 2994
rect 5460 2446 5488 3878
rect 5644 3126 5672 4082
rect 5724 3596 5776 3602
rect 5724 3538 5776 3544
rect 5632 3120 5684 3126
rect 5632 3062 5684 3068
rect 5736 3058 5764 3538
rect 5828 3534 5856 5510
rect 6092 5092 6144 5098
rect 6092 5034 6144 5040
rect 6104 4826 6132 5034
rect 6196 5030 6224 5714
rect 6748 5166 6776 6190
rect 6920 5704 6972 5710
rect 6920 5646 6972 5652
rect 7196 5704 7248 5710
rect 7300 5692 7328 7346
rect 7484 7274 7512 7346
rect 7472 7268 7524 7274
rect 7472 7210 7524 7216
rect 7380 6656 7432 6662
rect 7380 6598 7432 6604
rect 7248 5664 7328 5692
rect 7196 5646 7248 5652
rect 6828 5568 6880 5574
rect 6828 5510 6880 5516
rect 6840 5234 6868 5510
rect 6932 5370 6960 5646
rect 6920 5364 6972 5370
rect 6920 5306 6972 5312
rect 7300 5302 7328 5664
rect 7288 5296 7340 5302
rect 7288 5238 7340 5244
rect 6828 5228 6880 5234
rect 6828 5170 6880 5176
rect 6920 5228 6972 5234
rect 6920 5170 6972 5176
rect 6276 5160 6328 5166
rect 6736 5160 6788 5166
rect 6276 5102 6328 5108
rect 6656 5120 6736 5148
rect 6184 5024 6236 5030
rect 6184 4966 6236 4972
rect 6092 4820 6144 4826
rect 6092 4762 6144 4768
rect 6196 4282 6224 4966
rect 6288 4826 6316 5102
rect 6276 4820 6328 4826
rect 6276 4762 6328 4768
rect 6656 4282 6684 5120
rect 6736 5102 6788 5108
rect 6736 5024 6788 5030
rect 6736 4966 6788 4972
rect 6748 4690 6776 4966
rect 6736 4684 6788 4690
rect 6736 4626 6788 4632
rect 6184 4276 6236 4282
rect 6184 4218 6236 4224
rect 6644 4276 6696 4282
rect 6644 4218 6696 4224
rect 6368 4208 6420 4214
rect 6932 4162 6960 5170
rect 7392 4554 7420 6598
rect 7484 5846 7512 7210
rect 8220 6905 8248 7346
rect 8206 6896 8262 6905
rect 8206 6831 8262 6840
rect 8024 6316 8076 6322
rect 8024 6258 8076 6264
rect 7472 5840 7524 5846
rect 7472 5782 7524 5788
rect 7484 5574 7512 5782
rect 8036 5778 8064 6258
rect 8206 6216 8262 6225
rect 8206 6151 8208 6160
rect 8260 6151 8262 6160
rect 8208 6122 8260 6128
rect 8024 5772 8076 5778
rect 8024 5714 8076 5720
rect 7656 5704 7708 5710
rect 7656 5646 7708 5652
rect 7472 5568 7524 5574
rect 7472 5510 7524 5516
rect 7668 5098 7696 5646
rect 7656 5092 7708 5098
rect 7656 5034 7708 5040
rect 8036 4826 8064 5714
rect 8208 5704 8260 5710
rect 8208 5646 8260 5652
rect 8220 5545 8248 5646
rect 8206 5536 8262 5545
rect 8206 5471 8262 5480
rect 8208 5228 8260 5234
rect 8208 5170 8260 5176
rect 8220 4865 8248 5170
rect 8206 4856 8262 4865
rect 8024 4820 8076 4826
rect 8206 4791 8262 4800
rect 8024 4762 8076 4768
rect 7380 4548 7432 4554
rect 7380 4490 7432 4496
rect 6368 4150 6420 4156
rect 6000 4072 6052 4078
rect 6000 4014 6052 4020
rect 5816 3528 5868 3534
rect 5816 3470 5868 3476
rect 6012 3058 6040 4014
rect 6276 3936 6328 3942
rect 6276 3878 6328 3884
rect 5540 3052 5592 3058
rect 5540 2994 5592 3000
rect 5724 3052 5776 3058
rect 5724 2994 5776 3000
rect 6000 3052 6052 3058
rect 6000 2994 6052 3000
rect 5552 2650 5580 2994
rect 5632 2848 5684 2854
rect 5632 2790 5684 2796
rect 5724 2848 5776 2854
rect 5724 2790 5776 2796
rect 5908 2848 5960 2854
rect 5908 2790 5960 2796
rect 5540 2644 5592 2650
rect 5540 2586 5592 2592
rect 5644 2582 5672 2790
rect 5632 2576 5684 2582
rect 5632 2518 5684 2524
rect 5736 2514 5764 2790
rect 5724 2508 5776 2514
rect 5724 2450 5776 2456
rect 5448 2440 5500 2446
rect 5448 2382 5500 2388
rect 5632 2372 5684 2378
rect 5632 2314 5684 2320
rect 5644 2258 5672 2314
rect 5920 2310 5948 2790
rect 6012 2514 6040 2994
rect 6288 2990 6316 3878
rect 6276 2984 6328 2990
rect 6276 2926 6328 2932
rect 6380 2650 6408 4150
rect 6840 4134 6960 4162
rect 6736 3392 6788 3398
rect 6736 3334 6788 3340
rect 6748 3126 6776 3334
rect 6736 3120 6788 3126
rect 6736 3062 6788 3068
rect 6840 2774 6868 4134
rect 7196 4072 7248 4078
rect 7196 4014 7248 4020
rect 6656 2746 6868 2774
rect 6656 2650 6684 2746
rect 6368 2644 6420 2650
rect 6368 2586 6420 2592
rect 6644 2644 6696 2650
rect 6644 2586 6696 2592
rect 6552 2576 6604 2582
rect 6552 2518 6604 2524
rect 6000 2508 6052 2514
rect 6000 2450 6052 2456
rect 6564 2446 6592 2518
rect 6656 2446 6684 2586
rect 7208 2446 7236 4014
rect 7392 3534 7420 4490
rect 8116 4072 8168 4078
rect 8116 4014 8168 4020
rect 7380 3528 7432 3534
rect 7300 3476 7380 3482
rect 7300 3470 7432 3476
rect 7472 3528 7524 3534
rect 7472 3470 7524 3476
rect 7300 3454 7420 3470
rect 7300 3126 7328 3454
rect 7380 3392 7432 3398
rect 7380 3334 7432 3340
rect 7288 3120 7340 3126
rect 7288 3062 7340 3068
rect 6552 2440 6604 2446
rect 6552 2382 6604 2388
rect 6644 2440 6696 2446
rect 6644 2382 6696 2388
rect 7196 2440 7248 2446
rect 7196 2382 7248 2388
rect 7300 2310 7328 3062
rect 7392 2582 7420 3334
rect 7484 2650 7512 3470
rect 8128 3194 8156 4014
rect 8206 3496 8262 3505
rect 8206 3431 8262 3440
rect 8116 3188 8168 3194
rect 8116 3130 8168 3136
rect 7838 2816 7894 2825
rect 7838 2751 7894 2760
rect 7852 2650 7880 2751
rect 7472 2644 7524 2650
rect 7472 2586 7524 2592
rect 7840 2644 7892 2650
rect 7840 2586 7892 2592
rect 7380 2576 7432 2582
rect 7380 2518 7432 2524
rect 8220 2446 8248 3431
rect 8208 2440 8260 2446
rect 8208 2382 8260 2388
rect 5368 2230 5672 2258
rect 5908 2304 5960 2310
rect 5908 2246 5960 2252
rect 6460 2304 6512 2310
rect 6460 2246 6512 2252
rect 7288 2304 7340 2310
rect 7288 2246 7340 2252
rect 5368 2106 5396 2230
rect 5356 2100 5408 2106
rect 5356 2042 5408 2048
rect 5184 1278 5304 1306
rect 5184 800 5212 1278
rect 6472 800 6500 2246
rect 3238 0 3294 800
rect 4526 0 4582 800
rect 5170 0 5226 800
rect 6458 0 6514 800
<< via2 >>
rect 4220 9274 4276 9276
rect 4300 9274 4356 9276
rect 4380 9274 4436 9276
rect 4460 9274 4516 9276
rect 4220 9222 4266 9274
rect 4266 9222 4276 9274
rect 4300 9222 4330 9274
rect 4330 9222 4342 9274
rect 4342 9222 4356 9274
rect 4380 9222 4394 9274
rect 4394 9222 4406 9274
rect 4406 9222 4436 9274
rect 4460 9222 4470 9274
rect 4470 9222 4516 9274
rect 4220 9220 4276 9222
rect 4300 9220 4356 9222
rect 4380 9220 4436 9222
rect 4460 9220 4516 9222
rect 4880 8730 4936 8732
rect 4960 8730 5016 8732
rect 5040 8730 5096 8732
rect 5120 8730 5176 8732
rect 4880 8678 4926 8730
rect 4926 8678 4936 8730
rect 4960 8678 4990 8730
rect 4990 8678 5002 8730
rect 5002 8678 5016 8730
rect 5040 8678 5054 8730
rect 5054 8678 5066 8730
rect 5066 8678 5096 8730
rect 5120 8678 5130 8730
rect 5130 8678 5176 8730
rect 4880 8676 4936 8678
rect 4960 8676 5016 8678
rect 5040 8676 5096 8678
rect 5120 8676 5176 8678
rect 1398 8200 1454 8256
rect 846 7656 902 7712
rect 938 6840 994 6896
rect 4220 8186 4276 8188
rect 4300 8186 4356 8188
rect 4380 8186 4436 8188
rect 4460 8186 4516 8188
rect 4220 8134 4266 8186
rect 4266 8134 4276 8186
rect 4300 8134 4330 8186
rect 4330 8134 4342 8186
rect 4342 8134 4356 8186
rect 4380 8134 4394 8186
rect 4394 8134 4406 8186
rect 4406 8134 4436 8186
rect 4460 8134 4470 8186
rect 4470 8134 4516 8186
rect 4220 8132 4276 8134
rect 4300 8132 4356 8134
rect 4380 8132 4436 8134
rect 4460 8132 4516 8134
rect 846 6024 902 6080
rect 1674 5480 1730 5536
rect 846 4936 902 4992
rect 4880 7642 4936 7644
rect 4960 7642 5016 7644
rect 5040 7642 5096 7644
rect 5120 7642 5176 7644
rect 4880 7590 4926 7642
rect 4926 7590 4936 7642
rect 4960 7590 4990 7642
rect 4990 7590 5002 7642
rect 5002 7590 5016 7642
rect 5040 7590 5054 7642
rect 5054 7590 5066 7642
rect 5066 7590 5096 7642
rect 5120 7590 5130 7642
rect 5130 7590 5176 7642
rect 4880 7588 4936 7590
rect 4960 7588 5016 7590
rect 5040 7588 5096 7590
rect 5120 7588 5176 7590
rect 4220 7098 4276 7100
rect 4300 7098 4356 7100
rect 4380 7098 4436 7100
rect 4460 7098 4516 7100
rect 4220 7046 4266 7098
rect 4266 7046 4276 7098
rect 4300 7046 4330 7098
rect 4330 7046 4342 7098
rect 4342 7046 4356 7098
rect 4380 7046 4394 7098
rect 4394 7046 4406 7098
rect 4406 7046 4436 7098
rect 4460 7046 4470 7098
rect 4470 7046 4516 7098
rect 4220 7044 4276 7046
rect 4300 7044 4356 7046
rect 4380 7044 4436 7046
rect 4460 7044 4516 7046
rect 4880 6554 4936 6556
rect 4960 6554 5016 6556
rect 5040 6554 5096 6556
rect 5120 6554 5176 6556
rect 4880 6502 4926 6554
rect 4926 6502 4936 6554
rect 4960 6502 4990 6554
rect 4990 6502 5002 6554
rect 5002 6502 5016 6554
rect 5040 6502 5054 6554
rect 5054 6502 5066 6554
rect 5066 6502 5096 6554
rect 5120 6502 5130 6554
rect 5130 6502 5176 6554
rect 4880 6500 4936 6502
rect 4960 6500 5016 6502
rect 5040 6500 5096 6502
rect 5120 6500 5176 6502
rect 4220 6010 4276 6012
rect 4300 6010 4356 6012
rect 4380 6010 4436 6012
rect 4460 6010 4516 6012
rect 4220 5958 4266 6010
rect 4266 5958 4276 6010
rect 4300 5958 4330 6010
rect 4330 5958 4342 6010
rect 4342 5958 4356 6010
rect 4380 5958 4394 6010
rect 4394 5958 4406 6010
rect 4406 5958 4436 6010
rect 4460 5958 4470 6010
rect 4470 5958 4516 6010
rect 4220 5956 4276 5958
rect 4300 5956 4356 5958
rect 4380 5956 4436 5958
rect 4460 5956 4516 5958
rect 846 3612 848 3632
rect 848 3612 900 3632
rect 900 3612 902 3632
rect 846 3576 902 3612
rect 4220 4922 4276 4924
rect 4300 4922 4356 4924
rect 4380 4922 4436 4924
rect 4460 4922 4516 4924
rect 4220 4870 4266 4922
rect 4266 4870 4276 4922
rect 4300 4870 4330 4922
rect 4330 4870 4342 4922
rect 4342 4870 4356 4922
rect 4380 4870 4394 4922
rect 4394 4870 4406 4922
rect 4406 4870 4436 4922
rect 4460 4870 4470 4922
rect 4470 4870 4516 4922
rect 4220 4868 4276 4870
rect 4300 4868 4356 4870
rect 4380 4868 4436 4870
rect 4460 4868 4516 4870
rect 4880 5466 4936 5468
rect 4960 5466 5016 5468
rect 5040 5466 5096 5468
rect 5120 5466 5176 5468
rect 4880 5414 4926 5466
rect 4926 5414 4936 5466
rect 4960 5414 4990 5466
rect 4990 5414 5002 5466
rect 5002 5414 5016 5466
rect 5040 5414 5054 5466
rect 5054 5414 5066 5466
rect 5066 5414 5096 5466
rect 5120 5414 5130 5466
rect 5130 5414 5176 5466
rect 4880 5412 4936 5414
rect 4960 5412 5016 5414
rect 5040 5412 5096 5414
rect 5120 5412 5176 5414
rect 8206 7520 8262 7576
rect 4880 4378 4936 4380
rect 4960 4378 5016 4380
rect 5040 4378 5096 4380
rect 5120 4378 5176 4380
rect 4880 4326 4926 4378
rect 4926 4326 4936 4378
rect 4960 4326 4990 4378
rect 4990 4326 5002 4378
rect 5002 4326 5016 4378
rect 5040 4326 5054 4378
rect 5054 4326 5066 4378
rect 5066 4326 5096 4378
rect 5120 4326 5130 4378
rect 5130 4326 5176 4378
rect 4880 4324 4936 4326
rect 4960 4324 5016 4326
rect 5040 4324 5096 4326
rect 5120 4324 5176 4326
rect 4618 4120 4674 4176
rect 4220 3834 4276 3836
rect 4300 3834 4356 3836
rect 4380 3834 4436 3836
rect 4460 3834 4516 3836
rect 4220 3782 4266 3834
rect 4266 3782 4276 3834
rect 4300 3782 4330 3834
rect 4330 3782 4342 3834
rect 4342 3782 4356 3834
rect 4380 3782 4394 3834
rect 4394 3782 4406 3834
rect 4406 3782 4436 3834
rect 4460 3782 4470 3834
rect 4470 3782 4516 3834
rect 4220 3780 4276 3782
rect 4300 3780 4356 3782
rect 4380 3780 4436 3782
rect 4460 3780 4516 3782
rect 4880 3290 4936 3292
rect 4960 3290 5016 3292
rect 5040 3290 5096 3292
rect 5120 3290 5176 3292
rect 4880 3238 4926 3290
rect 4926 3238 4936 3290
rect 4960 3238 4990 3290
rect 4990 3238 5002 3290
rect 5002 3238 5016 3290
rect 5040 3238 5054 3290
rect 5054 3238 5066 3290
rect 5066 3238 5096 3290
rect 5120 3238 5130 3290
rect 5130 3238 5176 3290
rect 4880 3236 4936 3238
rect 4960 3236 5016 3238
rect 5040 3236 5096 3238
rect 5120 3236 5176 3238
rect 4220 2746 4276 2748
rect 4300 2746 4356 2748
rect 4380 2746 4436 2748
rect 4460 2746 4516 2748
rect 4220 2694 4266 2746
rect 4266 2694 4276 2746
rect 4300 2694 4330 2746
rect 4330 2694 4342 2746
rect 4342 2694 4356 2746
rect 4380 2694 4394 2746
rect 4394 2694 4406 2746
rect 4406 2694 4436 2746
rect 4460 2694 4470 2746
rect 4470 2694 4516 2746
rect 4220 2692 4276 2694
rect 4300 2692 4356 2694
rect 4380 2692 4436 2694
rect 4460 2692 4516 2694
rect 4880 2202 4936 2204
rect 4960 2202 5016 2204
rect 5040 2202 5096 2204
rect 5120 2202 5176 2204
rect 4880 2150 4926 2202
rect 4926 2150 4936 2202
rect 4960 2150 4990 2202
rect 4990 2150 5002 2202
rect 5002 2150 5016 2202
rect 5040 2150 5054 2202
rect 5054 2150 5066 2202
rect 5066 2150 5096 2202
rect 5120 2150 5130 2202
rect 5130 2150 5176 2202
rect 4880 2148 4936 2150
rect 4960 2148 5016 2150
rect 5040 2148 5096 2150
rect 5120 2148 5176 2150
rect 8206 6840 8262 6896
rect 8206 6180 8262 6216
rect 8206 6160 8208 6180
rect 8208 6160 8260 6180
rect 8260 6160 8262 6180
rect 8206 5480 8262 5536
rect 8206 4800 8262 4856
rect 8206 3440 8262 3496
rect 7838 2760 7894 2816
<< metal3 >>
rect 4210 9280 4526 9281
rect 4210 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4526 9280
rect 4210 9215 4526 9216
rect 4870 8736 5186 8737
rect 4870 8672 4876 8736
rect 4940 8672 4956 8736
rect 5020 8672 5036 8736
rect 5100 8672 5116 8736
rect 5180 8672 5186 8736
rect 4870 8671 5186 8672
rect 0 8258 800 8288
rect 1393 8258 1459 8261
rect 0 8256 1459 8258
rect 0 8200 1398 8256
rect 1454 8200 1459 8256
rect 0 8198 1459 8200
rect 0 8168 800 8198
rect 1393 8195 1459 8198
rect 4210 8192 4526 8193
rect 4210 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4526 8192
rect 4210 8127 4526 8128
rect 841 7714 907 7717
rect 798 7712 907 7714
rect 798 7656 846 7712
rect 902 7656 907 7712
rect 798 7651 907 7656
rect 798 7608 858 7651
rect 0 7518 858 7608
rect 4870 7648 5186 7649
rect 4870 7584 4876 7648
rect 4940 7584 4956 7648
rect 5020 7584 5036 7648
rect 5100 7584 5116 7648
rect 5180 7584 5186 7648
rect 4870 7583 5186 7584
rect 8201 7578 8267 7581
rect 8875 7578 9675 7608
rect 8201 7576 9675 7578
rect 8201 7520 8206 7576
rect 8262 7520 9675 7576
rect 8201 7518 9675 7520
rect 0 7488 800 7518
rect 8201 7515 8267 7518
rect 8875 7488 9675 7518
rect 4210 7104 4526 7105
rect 4210 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4526 7104
rect 4210 7039 4526 7040
rect 0 6898 800 6928
rect 933 6898 999 6901
rect 0 6896 999 6898
rect 0 6840 938 6896
rect 994 6840 999 6896
rect 0 6838 999 6840
rect 0 6808 800 6838
rect 933 6835 999 6838
rect 8201 6898 8267 6901
rect 8875 6898 9675 6928
rect 8201 6896 9675 6898
rect 8201 6840 8206 6896
rect 8262 6840 9675 6896
rect 8201 6838 9675 6840
rect 8201 6835 8267 6838
rect 8875 6808 9675 6838
rect 4870 6560 5186 6561
rect 4870 6496 4876 6560
rect 4940 6496 4956 6560
rect 5020 6496 5036 6560
rect 5100 6496 5116 6560
rect 5180 6496 5186 6560
rect 4870 6495 5186 6496
rect 0 6218 800 6248
rect 8201 6218 8267 6221
rect 8875 6218 9675 6248
rect 0 6128 858 6218
rect 8201 6216 9675 6218
rect 8201 6160 8206 6216
rect 8262 6160 9675 6216
rect 8201 6158 9675 6160
rect 8201 6155 8267 6158
rect 8875 6128 9675 6158
rect 798 6085 858 6128
rect 798 6080 907 6085
rect 798 6024 846 6080
rect 902 6024 907 6080
rect 798 6022 907 6024
rect 841 6019 907 6022
rect 4210 6016 4526 6017
rect 4210 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4526 6016
rect 4210 5951 4526 5952
rect 0 5538 800 5568
rect 1669 5538 1735 5541
rect 0 5536 1735 5538
rect 0 5480 1674 5536
rect 1730 5480 1735 5536
rect 0 5478 1735 5480
rect 0 5448 800 5478
rect 1669 5475 1735 5478
rect 8201 5538 8267 5541
rect 8875 5538 9675 5568
rect 8201 5536 9675 5538
rect 8201 5480 8206 5536
rect 8262 5480 9675 5536
rect 8201 5478 9675 5480
rect 8201 5475 8267 5478
rect 4870 5472 5186 5473
rect 4870 5408 4876 5472
rect 4940 5408 4956 5472
rect 5020 5408 5036 5472
rect 5100 5408 5116 5472
rect 5180 5408 5186 5472
rect 8875 5448 9675 5478
rect 4870 5407 5186 5408
rect 841 4994 907 4997
rect 798 4992 907 4994
rect 798 4936 846 4992
rect 902 4936 907 4992
rect 798 4931 907 4936
rect 798 4888 858 4931
rect 0 4798 858 4888
rect 4210 4928 4526 4929
rect 4210 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4526 4928
rect 4210 4863 4526 4864
rect 8201 4858 8267 4861
rect 8875 4858 9675 4888
rect 8201 4856 9675 4858
rect 8201 4800 8206 4856
rect 8262 4800 9675 4856
rect 8201 4798 9675 4800
rect 0 4768 800 4798
rect 8201 4795 8267 4798
rect 8875 4768 9675 4798
rect 4870 4384 5186 4385
rect 4870 4320 4876 4384
rect 4940 4320 4956 4384
rect 5020 4320 5036 4384
rect 5100 4320 5116 4384
rect 5180 4320 5186 4384
rect 4870 4319 5186 4320
rect 0 4178 800 4208
rect 4613 4178 4679 4181
rect 0 4176 4679 4178
rect 0 4120 4618 4176
rect 4674 4120 4679 4176
rect 0 4118 4679 4120
rect 0 4088 800 4118
rect 4613 4115 4679 4118
rect 4210 3840 4526 3841
rect 4210 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4526 3840
rect 4210 3775 4526 3776
rect 841 3634 907 3637
rect 798 3632 907 3634
rect 798 3576 846 3632
rect 902 3576 907 3632
rect 798 3571 907 3576
rect 798 3528 858 3571
rect 0 3438 858 3528
rect 8201 3498 8267 3501
rect 8875 3498 9675 3528
rect 8201 3496 9675 3498
rect 8201 3440 8206 3496
rect 8262 3440 9675 3496
rect 8201 3438 9675 3440
rect 0 3408 800 3438
rect 8201 3435 8267 3438
rect 8875 3408 9675 3438
rect 4870 3296 5186 3297
rect 4870 3232 4876 3296
rect 4940 3232 4956 3296
rect 5020 3232 5036 3296
rect 5100 3232 5116 3296
rect 5180 3232 5186 3296
rect 4870 3231 5186 3232
rect 7833 2818 7899 2821
rect 8875 2818 9675 2848
rect 7833 2816 9675 2818
rect 7833 2760 7838 2816
rect 7894 2760 9675 2816
rect 7833 2758 9675 2760
rect 7833 2755 7899 2758
rect 4210 2752 4526 2753
rect 4210 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4526 2752
rect 8875 2728 9675 2758
rect 4210 2687 4526 2688
rect 4870 2208 5186 2209
rect 4870 2144 4876 2208
rect 4940 2144 4956 2208
rect 5020 2144 5036 2208
rect 5100 2144 5116 2208
rect 5180 2144 5186 2208
rect 4870 2143 5186 2144
<< via3 >>
rect 4216 9276 4280 9280
rect 4216 9220 4220 9276
rect 4220 9220 4276 9276
rect 4276 9220 4280 9276
rect 4216 9216 4280 9220
rect 4296 9276 4360 9280
rect 4296 9220 4300 9276
rect 4300 9220 4356 9276
rect 4356 9220 4360 9276
rect 4296 9216 4360 9220
rect 4376 9276 4440 9280
rect 4376 9220 4380 9276
rect 4380 9220 4436 9276
rect 4436 9220 4440 9276
rect 4376 9216 4440 9220
rect 4456 9276 4520 9280
rect 4456 9220 4460 9276
rect 4460 9220 4516 9276
rect 4516 9220 4520 9276
rect 4456 9216 4520 9220
rect 4876 8732 4940 8736
rect 4876 8676 4880 8732
rect 4880 8676 4936 8732
rect 4936 8676 4940 8732
rect 4876 8672 4940 8676
rect 4956 8732 5020 8736
rect 4956 8676 4960 8732
rect 4960 8676 5016 8732
rect 5016 8676 5020 8732
rect 4956 8672 5020 8676
rect 5036 8732 5100 8736
rect 5036 8676 5040 8732
rect 5040 8676 5096 8732
rect 5096 8676 5100 8732
rect 5036 8672 5100 8676
rect 5116 8732 5180 8736
rect 5116 8676 5120 8732
rect 5120 8676 5176 8732
rect 5176 8676 5180 8732
rect 5116 8672 5180 8676
rect 4216 8188 4280 8192
rect 4216 8132 4220 8188
rect 4220 8132 4276 8188
rect 4276 8132 4280 8188
rect 4216 8128 4280 8132
rect 4296 8188 4360 8192
rect 4296 8132 4300 8188
rect 4300 8132 4356 8188
rect 4356 8132 4360 8188
rect 4296 8128 4360 8132
rect 4376 8188 4440 8192
rect 4376 8132 4380 8188
rect 4380 8132 4436 8188
rect 4436 8132 4440 8188
rect 4376 8128 4440 8132
rect 4456 8188 4520 8192
rect 4456 8132 4460 8188
rect 4460 8132 4516 8188
rect 4516 8132 4520 8188
rect 4456 8128 4520 8132
rect 4876 7644 4940 7648
rect 4876 7588 4880 7644
rect 4880 7588 4936 7644
rect 4936 7588 4940 7644
rect 4876 7584 4940 7588
rect 4956 7644 5020 7648
rect 4956 7588 4960 7644
rect 4960 7588 5016 7644
rect 5016 7588 5020 7644
rect 4956 7584 5020 7588
rect 5036 7644 5100 7648
rect 5036 7588 5040 7644
rect 5040 7588 5096 7644
rect 5096 7588 5100 7644
rect 5036 7584 5100 7588
rect 5116 7644 5180 7648
rect 5116 7588 5120 7644
rect 5120 7588 5176 7644
rect 5176 7588 5180 7644
rect 5116 7584 5180 7588
rect 4216 7100 4280 7104
rect 4216 7044 4220 7100
rect 4220 7044 4276 7100
rect 4276 7044 4280 7100
rect 4216 7040 4280 7044
rect 4296 7100 4360 7104
rect 4296 7044 4300 7100
rect 4300 7044 4356 7100
rect 4356 7044 4360 7100
rect 4296 7040 4360 7044
rect 4376 7100 4440 7104
rect 4376 7044 4380 7100
rect 4380 7044 4436 7100
rect 4436 7044 4440 7100
rect 4376 7040 4440 7044
rect 4456 7100 4520 7104
rect 4456 7044 4460 7100
rect 4460 7044 4516 7100
rect 4516 7044 4520 7100
rect 4456 7040 4520 7044
rect 4876 6556 4940 6560
rect 4876 6500 4880 6556
rect 4880 6500 4936 6556
rect 4936 6500 4940 6556
rect 4876 6496 4940 6500
rect 4956 6556 5020 6560
rect 4956 6500 4960 6556
rect 4960 6500 5016 6556
rect 5016 6500 5020 6556
rect 4956 6496 5020 6500
rect 5036 6556 5100 6560
rect 5036 6500 5040 6556
rect 5040 6500 5096 6556
rect 5096 6500 5100 6556
rect 5036 6496 5100 6500
rect 5116 6556 5180 6560
rect 5116 6500 5120 6556
rect 5120 6500 5176 6556
rect 5176 6500 5180 6556
rect 5116 6496 5180 6500
rect 4216 6012 4280 6016
rect 4216 5956 4220 6012
rect 4220 5956 4276 6012
rect 4276 5956 4280 6012
rect 4216 5952 4280 5956
rect 4296 6012 4360 6016
rect 4296 5956 4300 6012
rect 4300 5956 4356 6012
rect 4356 5956 4360 6012
rect 4296 5952 4360 5956
rect 4376 6012 4440 6016
rect 4376 5956 4380 6012
rect 4380 5956 4436 6012
rect 4436 5956 4440 6012
rect 4376 5952 4440 5956
rect 4456 6012 4520 6016
rect 4456 5956 4460 6012
rect 4460 5956 4516 6012
rect 4516 5956 4520 6012
rect 4456 5952 4520 5956
rect 4876 5468 4940 5472
rect 4876 5412 4880 5468
rect 4880 5412 4936 5468
rect 4936 5412 4940 5468
rect 4876 5408 4940 5412
rect 4956 5468 5020 5472
rect 4956 5412 4960 5468
rect 4960 5412 5016 5468
rect 5016 5412 5020 5468
rect 4956 5408 5020 5412
rect 5036 5468 5100 5472
rect 5036 5412 5040 5468
rect 5040 5412 5096 5468
rect 5096 5412 5100 5468
rect 5036 5408 5100 5412
rect 5116 5468 5180 5472
rect 5116 5412 5120 5468
rect 5120 5412 5176 5468
rect 5176 5412 5180 5468
rect 5116 5408 5180 5412
rect 4216 4924 4280 4928
rect 4216 4868 4220 4924
rect 4220 4868 4276 4924
rect 4276 4868 4280 4924
rect 4216 4864 4280 4868
rect 4296 4924 4360 4928
rect 4296 4868 4300 4924
rect 4300 4868 4356 4924
rect 4356 4868 4360 4924
rect 4296 4864 4360 4868
rect 4376 4924 4440 4928
rect 4376 4868 4380 4924
rect 4380 4868 4436 4924
rect 4436 4868 4440 4924
rect 4376 4864 4440 4868
rect 4456 4924 4520 4928
rect 4456 4868 4460 4924
rect 4460 4868 4516 4924
rect 4516 4868 4520 4924
rect 4456 4864 4520 4868
rect 4876 4380 4940 4384
rect 4876 4324 4880 4380
rect 4880 4324 4936 4380
rect 4936 4324 4940 4380
rect 4876 4320 4940 4324
rect 4956 4380 5020 4384
rect 4956 4324 4960 4380
rect 4960 4324 5016 4380
rect 5016 4324 5020 4380
rect 4956 4320 5020 4324
rect 5036 4380 5100 4384
rect 5036 4324 5040 4380
rect 5040 4324 5096 4380
rect 5096 4324 5100 4380
rect 5036 4320 5100 4324
rect 5116 4380 5180 4384
rect 5116 4324 5120 4380
rect 5120 4324 5176 4380
rect 5176 4324 5180 4380
rect 5116 4320 5180 4324
rect 4216 3836 4280 3840
rect 4216 3780 4220 3836
rect 4220 3780 4276 3836
rect 4276 3780 4280 3836
rect 4216 3776 4280 3780
rect 4296 3836 4360 3840
rect 4296 3780 4300 3836
rect 4300 3780 4356 3836
rect 4356 3780 4360 3836
rect 4296 3776 4360 3780
rect 4376 3836 4440 3840
rect 4376 3780 4380 3836
rect 4380 3780 4436 3836
rect 4436 3780 4440 3836
rect 4376 3776 4440 3780
rect 4456 3836 4520 3840
rect 4456 3780 4460 3836
rect 4460 3780 4516 3836
rect 4516 3780 4520 3836
rect 4456 3776 4520 3780
rect 4876 3292 4940 3296
rect 4876 3236 4880 3292
rect 4880 3236 4936 3292
rect 4936 3236 4940 3292
rect 4876 3232 4940 3236
rect 4956 3292 5020 3296
rect 4956 3236 4960 3292
rect 4960 3236 5016 3292
rect 5016 3236 5020 3292
rect 4956 3232 5020 3236
rect 5036 3292 5100 3296
rect 5036 3236 5040 3292
rect 5040 3236 5096 3292
rect 5096 3236 5100 3292
rect 5036 3232 5100 3236
rect 5116 3292 5180 3296
rect 5116 3236 5120 3292
rect 5120 3236 5176 3292
rect 5176 3236 5180 3292
rect 5116 3232 5180 3236
rect 4216 2748 4280 2752
rect 4216 2692 4220 2748
rect 4220 2692 4276 2748
rect 4276 2692 4280 2748
rect 4216 2688 4280 2692
rect 4296 2748 4360 2752
rect 4296 2692 4300 2748
rect 4300 2692 4356 2748
rect 4356 2692 4360 2748
rect 4296 2688 4360 2692
rect 4376 2748 4440 2752
rect 4376 2692 4380 2748
rect 4380 2692 4436 2748
rect 4436 2692 4440 2748
rect 4376 2688 4440 2692
rect 4456 2748 4520 2752
rect 4456 2692 4460 2748
rect 4460 2692 4516 2748
rect 4516 2692 4520 2748
rect 4456 2688 4520 2692
rect 4876 2204 4940 2208
rect 4876 2148 4880 2204
rect 4880 2148 4936 2204
rect 4936 2148 4940 2204
rect 4876 2144 4940 2148
rect 4956 2204 5020 2208
rect 4956 2148 4960 2204
rect 4960 2148 5016 2204
rect 5016 2148 5020 2204
rect 4956 2144 5020 2148
rect 5036 2204 5100 2208
rect 5036 2148 5040 2204
rect 5040 2148 5096 2204
rect 5096 2148 5100 2204
rect 5036 2144 5100 2148
rect 5116 2204 5180 2208
rect 5116 2148 5120 2204
rect 5120 2148 5176 2204
rect 5176 2148 5180 2204
rect 5116 2144 5180 2148
<< metal4 >>
rect 4208 9280 4528 9296
rect 4208 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4528 9280
rect 4208 8192 4528 9216
rect 4208 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4528 8192
rect 4208 7104 4528 8128
rect 4208 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4528 7104
rect 4208 6016 4528 7040
rect 4208 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4528 6016
rect 4208 4928 4528 5952
rect 4208 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4528 4928
rect 4208 3840 4528 4864
rect 4208 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4528 3840
rect 4208 2752 4528 3776
rect 4208 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4528 2752
rect 4208 2128 4528 2688
rect 4868 8736 5188 9296
rect 4868 8672 4876 8736
rect 4940 8672 4956 8736
rect 5020 8672 5036 8736
rect 5100 8672 5116 8736
rect 5180 8672 5188 8736
rect 4868 7648 5188 8672
rect 4868 7584 4876 7648
rect 4940 7584 4956 7648
rect 5020 7584 5036 7648
rect 5100 7584 5116 7648
rect 5180 7584 5188 7648
rect 4868 6560 5188 7584
rect 4868 6496 4876 6560
rect 4940 6496 4956 6560
rect 5020 6496 5036 6560
rect 5100 6496 5116 6560
rect 5180 6496 5188 6560
rect 4868 5472 5188 6496
rect 4868 5408 4876 5472
rect 4940 5408 4956 5472
rect 5020 5408 5036 5472
rect 5100 5408 5116 5472
rect 5180 5408 5188 5472
rect 4868 4384 5188 5408
rect 4868 4320 4876 4384
rect 4940 4320 4956 4384
rect 5020 4320 5036 4384
rect 5100 4320 5116 4384
rect 5180 4320 5188 4384
rect 4868 3296 5188 4320
rect 4868 3232 4876 3296
rect 4940 3232 4956 3296
rect 5020 3232 5036 3296
rect 5100 3232 5116 3296
rect 5180 3232 5188 3296
rect 4868 2208 5188 3232
rect 4868 2144 4876 2208
rect 4940 2144 4956 2208
rect 5020 2144 5036 2208
rect 5100 2144 5116 2208
rect 5180 2144 5188 2208
rect 4868 2128 5188 2144
use sky130_fd_sc_hd__inv_2  _054_
timestamp 0
transform -1 0 7268 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _055_
timestamp 0
transform -1 0 7544 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _056_
timestamp 0
transform 1 0 2024 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_2  _057_
timestamp 0
transform 1 0 7360 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__and2b_2  _058_
timestamp 0
transform -1 0 7636 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _059_
timestamp 0
transform -1 0 6992 0 1 2176
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _060_
timestamp 0
transform 1 0 6348 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__nand2b_1  _061_
timestamp 0
transform 1 0 4048 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _062_
timestamp 0
transform 1 0 4508 0 1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _063_
timestamp 0
transform 1 0 5796 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _064_
timestamp 0
transform -1 0 5428 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _065_
timestamp 0
transform 1 0 5152 0 -1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _066_
timestamp 0
transform 1 0 4968 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _067_
timestamp 0
transform 1 0 4324 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__xor2_1  _068_
timestamp 0
transform 1 0 1380 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _069_
timestamp 0
transform -1 0 3864 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _070_
timestamp 0
transform -1 0 3588 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _071_
timestamp 0
transform 1 0 2576 0 1 2176
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _072_
timestamp 0
transform 1 0 2668 0 1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _073_
timestamp 0
transform 1 0 1380 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _074_
timestamp 0
transform 1 0 4048 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _075_
timestamp 0
transform 1 0 2116 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _076_
timestamp 0
transform 1 0 2392 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _077_
timestamp 0
transform 1 0 2024 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__a221o_1  _078_
timestamp 0
transform 1 0 2024 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__o21bai_1  _079_
timestamp 0
transform -1 0 4048 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__o31ai_2  _080_
timestamp 0
transform -1 0 4692 0 1 4352
box -38 -48 958 592
use sky130_fd_sc_hd__and2b_1  _081_
timestamp 0
transform -1 0 6256 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _082_
timestamp 0
transform -1 0 5704 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _083_
timestamp 0
transform -1 0 5152 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _084_
timestamp 0
transform 1 0 5704 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _085_
timestamp 0
transform 1 0 6164 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _086_
timestamp 0
transform -1 0 7360 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _087_
timestamp 0
transform 1 0 6348 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _088_
timestamp 0
transform 1 0 5704 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _089_
timestamp 0
transform -1 0 5704 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _090_
timestamp 0
transform 1 0 5704 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _091_
timestamp 0
transform 1 0 5980 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _092_
timestamp 0
transform -1 0 7636 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _093_
timestamp 0
transform 1 0 6624 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _094_
timestamp 0
transform 1 0 4416 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _095_
timestamp 0
transform 1 0 4968 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _096_
timestamp 0
transform -1 0 5796 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__o21ba_1  _097_
timestamp 0
transform 1 0 5520 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _098_
timestamp 0
transform 1 0 4876 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _099_
timestamp 0
transform -1 0 5612 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _100_
timestamp 0
transform 1 0 6348 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _101_
timestamp 0
transform -1 0 5336 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _102_
timestamp 0
transform 1 0 4048 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _103_
timestamp 0
transform 1 0 4048 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _104_
timestamp 0
transform 1 0 1840 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _105_
timestamp 0
transform -1 0 3312 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _106_
timestamp 0
transform 1 0 2024 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _107_
timestamp 0
transform 1 0 2484 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__dfrtp_1  _108_
timestamp 0
transform 1 0 6440 0 -1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _109_
timestamp 0
transform -1 0 5152 0 -1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _110_
timestamp 0
transform -1 0 3312 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _111_
timestamp 0
transform 1 0 2484 0 -1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _112_
timestamp 0
transform 1 0 6440 0 1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _113_
timestamp 0
transform 1 0 6440 0 1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _114_
timestamp 0
transform 1 0 3772 0 1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _115_
timestamp 0
transform -1 0 3220 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_clk
timestamp 0
transform 1 0 4508 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f_clk
timestamp 0
transform 1 0 5428 0 1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f_clk
timestamp 0
transform -1 0 5704 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_4  clkload0
timestamp 0
transform 1 0 5428 0 -1 4352
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_3
timestamp 0
transform 1 0 1380 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_15
timestamp 0
transform 1 0 2484 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_23
timestamp 0
transform 1 0 3220 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_27
timestamp 0
transform 1 0 3588 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_29
timestamp 0
transform 1 0 3772 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_37
timestamp 0
transform 1 0 4508 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_41
timestamp 0
transform 1 0 4876 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_51
timestamp 0
transform 1 0 5796 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_55
timestamp 0
transform 1 0 6164 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_70
timestamp 0
transform 1 0 7544 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_54
timestamp 0
transform 1 0 6072 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_57
timestamp 0
transform 1 0 6348 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2_6
timestamp 0
transform 1 0 1656 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_14
timestamp 0
transform 1 0 2392 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_24
timestamp 0
transform 1 0 3312 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_29
timestamp 0
transform 1 0 3772 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_44
timestamp 0
transform 1 0 5152 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2_70
timestamp 0
transform 1 0 7544 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3_13
timestamp 0
transform 1 0 2300 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_21
timestamp 0
transform 1 0 3036 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_30
timestamp 0
transform 1 0 3864 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_34
timestamp 0
transform 1 0 4232 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_53
timestamp 0
transform 1 0 5980 0 -1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_61
timestamp 0
transform 1 0 6716 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_73
timestamp 0
transform 1 0 7820 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_77
timestamp 0
transform 1 0 8188 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4_3
timestamp 0
transform 1 0 1380 0 1 4352
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_15
timestamp 0
transform 1 0 2484 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_27
timestamp 0
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4_39
timestamp 0
transform 1 0 4692 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_43
timestamp 0
transform 1 0 5060 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_7
timestamp 0
transform 1 0 1748 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_18
timestamp 0
transform 1 0 2760 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_35
timestamp 0
transform 1 0 4324 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_71
timestamp 0
transform 1 0 7636 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_6_18
timestamp 0
transform 1 0 2760 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_26
timestamp 0
transform 1 0 3496 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_6_29
timestamp 0
transform 1 0 3772 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_57
timestamp 0
transform 1 0 6348 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_73
timestamp 0
transform 1 0 7820 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_9
timestamp 0
transform 1 0 1932 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_35
timestamp 0
transform 1 0 4324 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_57
timestamp 0
transform 1 0 6348 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_67
timestamp 0
transform 1 0 7268 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_9
timestamp 0
transform 1 0 1932 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_8_17
timestamp 0
transform 1 0 2668 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_25
timestamp 0
transform 1 0 3404 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_49
timestamp 0
transform 1 0 5612 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_23
timestamp 0
transform 1 0 3220 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_29
timestamp 0
transform 1 0 3772 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_50
timestamp 0
transform 1 0 5704 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_57
timestamp 0
transform 1 0 6348 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_63
timestamp 0
transform 1 0 6900 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_71
timestamp 0
transform 1 0 7636 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_10_6
timestamp 0
transform 1 0 1656 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_14
timestamp 0
transform 1 0 2392 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_21
timestamp 0
transform 1 0 3036 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_27
timestamp 0
transform 1 0 3588 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_29
timestamp 0
transform 1 0 3772 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_49
timestamp 0
transform 1 0 5612 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_62
timestamp 0
transform 1 0 6808 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_74
timestamp 0
transform 1 0 7912 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_6
timestamp 0
transform 1 0 1656 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_15
timestamp 0
transform 1 0 2484 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_11_24
timestamp 0
transform 1 0 3312 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_51
timestamp 0
transform 1 0 5796 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_55
timestamp 0
transform 1 0 6164 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_57
timestamp 0
transform 1 0 6348 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_11_69
timestamp 0
transform 1 0 7452 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_77
timestamp 0
transform 1 0 8188 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_3
timestamp 0
transform 1 0 1380 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_15
timestamp 0
transform 1 0 2484 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_27
timestamp 0
transform 1 0 3588 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_29
timestamp 0
transform 1 0 3772 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_37
timestamp 0
transform 1 0 4508 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_41
timestamp 0
transform 1 0 4876 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_48
timestamp 0
transform 1 0 5520 0 1 8704
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_57
timestamp 0
transform 1 0 6348 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_69
timestamp 0
transform 1 0 7452 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_77
timestamp 0
transform 1 0 8188 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input1
timestamp 0
transform -1 0 7544 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input2
timestamp 0
transform -1 0 5796 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input3
timestamp 0
transform 1 0 3312 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input4
timestamp 0
transform -1 0 1656 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input5
timestamp 0
transform 1 0 8004 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input6
timestamp 0
transform 1 0 8004 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input7
timestamp 0
transform 1 0 5244 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input8
timestamp 0
transform -1 0 1656 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input9
timestamp 0
transform -1 0 8280 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input10
timestamp 0
transform 1 0 1380 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input11
timestamp 0
transform -1 0 8280 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input12
timestamp 0
transform 1 0 1380 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__buf_1  output13
timestamp 0
transform 1 0 7636 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  output14
timestamp 0
transform -1 0 4876 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  output15
timestamp 0
transform -1 0 1656 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  output16
timestamp 0
transform -1 0 1932 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  output17
timestamp 0
transform 1 0 8004 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  output18
timestamp 0
transform 1 0 8004 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  output19
timestamp 0
transform -1 0 4876 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  output20
timestamp 0
transform -1 0 1656 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Left_13
timestamp 0
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Right_0
timestamp 0
transform -1 0 8556 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Left_14
timestamp 0
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Right_1
timestamp 0
transform -1 0 8556 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Left_15
timestamp 0
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Right_2
timestamp 0
transform -1 0 8556 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Left_16
timestamp 0
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Right_3
timestamp 0
transform -1 0 8556 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Left_17
timestamp 0
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Right_4
timestamp 0
transform -1 0 8556 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Left_18
timestamp 0
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Right_5
timestamp 0
transform -1 0 8556 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Left_19
timestamp 0
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Right_6
timestamp 0
transform -1 0 8556 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Left_20
timestamp 0
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Right_7
timestamp 0
transform -1 0 8556 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Left_21
timestamp 0
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Right_8
timestamp 0
transform -1 0 8556 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Left_22
timestamp 0
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Right_9
timestamp 0
transform -1 0 8556 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Left_23
timestamp 0
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Right_10
timestamp 0
transform -1 0 8556 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Left_24
timestamp 0
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Right_11
timestamp 0
transform -1 0 8556 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Left_25
timestamp 0
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Right_12
timestamp 0
transform -1 0 8556 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_26
timestamp 0
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_27
timestamp 0
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_28
timestamp 0
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_29
timestamp 0
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_30
timestamp 0
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_31
timestamp 0
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_32
timestamp 0
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_33
timestamp 0
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_34
timestamp 0
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_35
timestamp 0
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_36
timestamp 0
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_37
timestamp 0
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_38
timestamp 0
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_39
timestamp 0
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_40
timestamp 0
transform 1 0 6256 0 1 8704
box -38 -48 130 592
<< labels >>
rlabel metal1 s 4830 8704 4830 8704 4 VGND
rlabel metal1 s 4830 9248 4830 9248 4 VPWR
rlabel metal1 s 6532 2958 6532 2958 4 _000_
rlabel metal1 s 4922 2618 4922 2618 4 _001_
rlabel metal2 s 2990 3230 2990 3230 4 _002_
rlabel metal2 s 2806 6052 2806 6052 4 _003_
rlabel metal2 s 6762 4828 6762 4828 4 _004_
rlabel metal1 s 6716 6426 6716 6426 4 _005_
rlabel metal1 s 3992 6970 3992 6970 4 _006_
rlabel metal2 s 2806 7582 2806 7582 4 _007_
rlabel metal1 s 6946 2448 6946 2448 4 _008_
rlabel metal1 s 6992 2550 6992 2550 4 _009_
rlabel metal1 s 2208 4250 2208 4250 4 _010_
rlabel metal1 s 2346 5576 2346 5576 4 _011_
rlabel metal2 s 4462 7854 4462 7854 4 _012_
rlabel metal2 s 6394 3400 6394 3400 4 _013_
rlabel metal1 s 4554 3638 4554 3638 4 _014_
rlabel metal1 s 5428 3570 5428 3570 4 _015_
rlabel metal1 s 5658 2278 5658 2278 4 _016_
rlabel metal1 s 5428 3910 5428 3910 4 _017_
rlabel metal1 s 5290 2414 5290 2414 4 _018_
rlabel metal2 s 4370 4420 4370 4420 4 _019_
rlabel metal1 s 3542 4080 3542 4080 4 _020_
rlabel metal1 s 3358 3570 3358 3570 4 _021_
rlabel metal2 s 3174 4386 3174 4386 4 _022_
rlabel metal2 s 3174 3060 3174 3060 4 _023_
rlabel metal2 s 1978 5440 1978 5440 4 _024_
rlabel metal2 s 4094 4794 4094 4794 4 _025_
rlabel metal1 s 2438 5134 2438 5134 4 _026_
rlabel metal1 s 2392 5270 2392 5270 4 _027_
rlabel metal2 s 2070 5372 2070 5372 4 _028_
rlabel metal2 s 3818 4794 3818 4794 4 _029_
rlabel metal1 s 5106 5338 5106 5338 4 _030_
rlabel metal1 s 5474 5168 5474 5168 4 _031_
rlabel metal1 s 5152 4794 5152 4794 4 _032_
rlabel metal2 s 5244 5202 5244 5202 4 _033_
rlabel metal2 s 6118 4930 6118 4930 4 _034_
rlabel metal2 s 6302 4964 6302 4964 4 _035_
rlabel metal2 s 6854 5372 6854 5372 4 _036_
rlabel metal1 s 6256 6766 6256 6766 4 _037_
rlabel metal2 s 5750 6052 5750 6052 4 _038_
rlabel metal1 s 6946 6324 6946 6324 4 _039_
rlabel metal2 s 6854 6460 6854 6460 4 _040_
rlabel metal2 s 7130 6732 7130 6732 4 _041_
rlabel metal1 s 4738 8398 4738 8398 4 _042_
rlabel metal1 s 5750 8432 5750 8432 4 _043_
rlabel metal1 s 4968 8602 4968 8602 4 _044_
rlabel metal1 s 5474 6222 5474 6222 4 _045_
rlabel metal1 s 5520 7854 5520 7854 4 _046_
rlabel metal2 s 4370 7820 4370 7820 4 _047_
rlabel metal1 s 4278 7990 4278 7990 4 _048_
rlabel metal1 s 4554 7956 4554 7956 4 _049_
rlabel metal1 s 3082 8432 3082 8432 4 _050_
rlabel metal1 s 2438 8364 2438 8364 4 _051_
rlabel metal2 s 2806 8058 2806 8058 4 _052_
rlabel metal1 s 2668 6970 2668 6970 4 _053_
rlabel metal2 s 4646 4879 4646 4879 4 clk
rlabel metal2 s 5842 4522 5842 4522 4 clknet_0_clk
rlabel metal1 s 5106 3094 5106 3094 4 clknet_1_0__leaf_clk
rlabel metal1 s 2530 6358 2530 6358 4 clknet_1_1__leaf_clk
rlabel metal3 s 8380 2788 8380 2788 4 count[0]
rlabel metal2 s 4554 1520 4554 1520 4 count[1]
rlabel metal3 s 0 3408 800 3528 4 count[2]
port 6 nsew
rlabel metal3 s 1188 5508 1188 5508 4 count[3]
rlabel metal3 s 8234 6171 8234 6171 4 count[4]
rlabel metal2 s 8234 7633 8234 7633 4 count[5]
rlabel metal2 s 4646 9571 4646 9571 4 count[6]
rlabel metal3 s 1050 8228 1050 8228 4 count[7]
rlabel metal2 s 6486 1520 6486 1520 4 data[0]
rlabel metal2 s 5198 1027 5198 1027 4 data[1]
rlabel metal2 s 3266 1622 3266 1622 4 data[2]
rlabel metal3 s 0 6128 800 6248 4 data[3]
port 15 nsew
rlabel metal2 s 8234 5015 8234 5015 4 data[4]
rlabel metal2 s 8234 7123 8234 7123 4 data[5]
rlabel metal1 s 5336 8942 5336 8942 4 data[6]
rlabel metal3 s 0 7488 800 7608 4 data[7]
port 19 nsew
rlabel metal2 s 8234 5593 8234 5593 4 enable
rlabel metal2 s 7498 3060 7498 3060 4 net1
rlabel metal1 s 1610 5100 1610 5100 4 net10
rlabel metal2 s 2530 3264 2530 3264 4 net11
rlabel metal1 s 1932 6970 1932 6970 4 net12
rlabel metal1 s 7682 2448 7682 2448 4 net13
rlabel metal1 s 5060 2482 5060 2482 4 net14
rlabel metal1 s 2392 4114 2392 4114 4 net15
rlabel metal2 s 1886 6018 1886 6018 4 net16
rlabel metal2 s 8050 5542 8050 5542 4 net17
rlabel metal2 s 6026 7106 6026 7106 4 net18
rlabel metal1 s 5290 7820 5290 7820 4 net19
rlabel metal1 s 5658 2618 5658 2618 4 net2
rlabel metal1 s 1840 6766 1840 6766 4 net20
rlabel metal1 s 3082 2414 3082 2414 4 net3
rlabel metal2 s 2532 5678 2532 5678 4 net4
rlabel metal1 s 7498 5338 7498 5338 4 net5
rlabel metal1 s 7222 7412 7222 7412 4 net6
rlabel metal1 s 4922 7922 4922 7922 4 net7
rlabel metal1 s 2024 7718 2024 7718 4 net8
rlabel metal1 s 7866 5678 7866 5678 4 net9
rlabel metal3 s 0 4768 800 4888 4 preload
port 21 nsew
rlabel metal3 s 8564 3468 8564 3468 4 resetn
rlabel metal1 s 1242 6766 1242 6766 4 up_down
flabel metal4 s 4868 2128 5188 9296 0 FreeSans 2400 90 0 0 VGND
port 1 nsew
flabel metal4 s 4208 2128 4528 9296 0 FreeSans 2400 90 0 0 VPWR
port 2 nsew
flabel metal3 s 0 4088 800 4208 0 FreeSans 600 0 0 0 clk
port 3 nsew
flabel metal3 s 8875 2728 9675 2848 0 FreeSans 600 0 0 0 count[0]
port 4 nsew
flabel metal2 s 4526 0 4582 800 0 FreeSans 280 90 0 0 count[1]
port 5 nsew
flabel metal3 s 400 3468 400 3468 0 FreeSans 600 0 0 0 count[2]
flabel metal3 s 0 5448 800 5568 0 FreeSans 600 0 0 0 count[3]
port 7 nsew
flabel metal3 s 8875 6128 9675 6248 0 FreeSans 600 0 0 0 count[4]
port 8 nsew
flabel metal3 s 8875 7488 9675 7608 0 FreeSans 600 0 0 0 count[5]
port 9 nsew
flabel metal2 s 4526 11019 4582 11819 0 FreeSans 280 90 0 0 count[6]
port 10 nsew
flabel metal3 s 0 8168 800 8288 0 FreeSans 600 0 0 0 count[7]
port 11 nsew
flabel metal2 s 6458 0 6514 800 0 FreeSans 280 90 0 0 data[0]
port 12 nsew
flabel metal2 s 5170 0 5226 800 0 FreeSans 280 90 0 0 data[1]
port 13 nsew
flabel metal2 s 3238 0 3294 800 0 FreeSans 280 90 0 0 data[2]
port 14 nsew
flabel metal3 s 400 6188 400 6188 0 FreeSans 600 0 0 0 data[3]
flabel metal3 s 8875 4768 9675 4888 0 FreeSans 600 0 0 0 data[4]
port 16 nsew
flabel metal3 s 8875 6808 9675 6928 0 FreeSans 600 0 0 0 data[5]
port 17 nsew
flabel metal2 s 5170 11019 5226 11819 0 FreeSans 280 90 0 0 data[6]
port 18 nsew
flabel metal3 s 400 7548 400 7548 0 FreeSans 600 0 0 0 data[7]
flabel metal3 s 8875 5448 9675 5568 0 FreeSans 600 0 0 0 enable
port 20 nsew
flabel metal3 s 400 4828 400 4828 0 FreeSans 600 0 0 0 preload
flabel metal3 s 8875 3408 9675 3528 0 FreeSans 600 0 0 0 resetn
port 22 nsew
flabel metal3 s 0 6808 800 6928 0 FreeSans 600 0 0 0 up_down
port 23 nsew
<< properties >>
string FIXED_BBOX 0 0 9675 11819
<< end >>
