* NGSPICE file created from counter.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_1 abstract view
.subckt sky130_fd_sc_hd__xor2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_1 abstract view
.subckt sky130_fd_sc_hd__dfrtp_1 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_1 abstract view
.subckt sky130_fd_sc_hd__buf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_1 abstract view
.subckt sky130_fd_sc_hd__nand2b_1 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_1 abstract view
.subckt sky130_fd_sc_hd__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_2 abstract view
.subckt sky130_fd_sc_hd__dfrtp_2 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_1 abstract view
.subckt sky130_fd_sc_hd__a31o_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_1 abstract view
.subckt sky130_fd_sc_hd__o21ba_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_1 abstract view
.subckt sky130_fd_sc_hd__o21bai_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VPWR VGND VPB VNB
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_1 abstract view
.subckt sky130_fd_sc_hd__and2b_1 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_1 abstract view
.subckt sky130_fd_sc_hd__a221o_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_1 abstract view
.subckt sky130_fd_sc_hd__o21ai_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_1 abstract view
.subckt sky130_fd_sc_hd__a22o_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_2 abstract view
.subckt sky130_fd_sc_hd__and2b_2 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_1 abstract view
.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_2 abstract view
.subckt sky130_fd_sc_hd__nor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_1 abstract view
.subckt sky130_fd_sc_hd__xnor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_1 abstract view
.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_1 abstract view
.subckt sky130_fd_sc_hd__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_2 abstract view
.subckt sky130_fd_sc_hd__o31ai_2 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

.subckt counter VGND VPWR clk count[0] count[1] count[2] count[3] count[4] count[5]
+ count[6] count[7] data[0] data[1] data[2] data[3] data[4] data[5] data[6] data[7]
+ enable preload resetn up_down
XFILLER_0_10_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_062_ net14 net12 VGND VGND VPWR VPWR _015_ sky130_fd_sc_hd__xor2_1
XPHY_EDGE_ROW_12_Left_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_114_ clknet_1_1__leaf_clk _006_ net11 VGND VGND VPWR VPWR net19 sky130_fd_sc_hd__dfrtp_1
Xoutput20 net20 VGND VGND VPWR VPWR count[7] sky130_fd_sc_hd__buf_1
XPHY_EDGE_ROW_12_Right_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_0_Left_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_113_ clknet_1_1__leaf_clk _005_ net11 VGND VGND VPWR VPWR net18 sky130_fd_sc_hd__dfrtp_1
X_061_ net12 net14 VGND VGND VPWR VPWR _014_ sky130_fd_sc_hd__nand2b_1
XPHY_EDGE_ROW_6_Right_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_6_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_6_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_11_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_10_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_9_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_8_35 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_060_ net13 _012_ _013_ VGND VGND VPWR VPWR _000_ sky130_fd_sc_hd__a21oi_1
X_112_ clknet_1_0__leaf_clk _004_ net11 VGND VGND VPWR VPWR net17 sky130_fd_sc_hd__dfrtp_1
X_111_ clknet_1_1__leaf_clk _003_ net11 VGND VGND VPWR VPWR net16 sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_4_Left_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_7_Left_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_110_ clknet_1_0__leaf_clk _002_ net11 VGND VGND VPWR VPWR net15 sky130_fd_sc_hd__dfrtp_2
XFILLER_0_1_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkload0 clknet_1_0__leaf_clk VGND VGND VPWR VPWR clkload0/X sky130_fd_sc_hd__clkbuf_4
Xoutput13 net13 VGND VGND VPWR VPWR count[0] sky130_fd_sc_hd__buf_1
XFILLER_0_4_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput14 net14 VGND VGND VPWR VPWR count[1] sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_2_29 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_099_ _044_ _046_ VGND VGND VPWR VPWR _047_ sky130_fd_sc_hd__nand2_1
XPHY_EDGE_ROW_1_Right_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput15 net15 VGND VGND VPWR VPWR count[2] sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_12_39 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_098_ _030_ _033_ _037_ _045_ VGND VGND VPWR VPWR _046_ sky130_fd_sc_hd__a31o_1
XFILLER_0_1_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_0_clk clk VGND VGND VPWR VPWR clknet_0_clk sky130_fd_sc_hd__clkbuf_16
Xoutput16 net16 VGND VGND VPWR VPWR count[3] sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_3_30 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_097_ net17 net18 net12 VGND VGND VPWR VPWR _045_ sky130_fd_sc_hd__o21ba_1
XPHY_EDGE_ROW_11_Left_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput17 net17 VGND VGND VPWR VPWR count[4] sky130_fd_sc_hd__buf_1
XFILLER_0_7_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_7_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_096_ _042_ _043_ VGND VGND VPWR VPWR _044_ sky130_fd_sc_hd__nor2_1
Xoutput18 net18 VGND VGND VPWR VPWR count[5] sky130_fd_sc_hd__buf_1
XPHY_EDGE_ROW_5_Right_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_079_ net15 net16 net12 VGND VGND VPWR VPWR _029_ sky130_fd_sc_hd__o21bai_1
XFILLER_0_4_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_095_ net19 net12 VGND VGND VPWR VPWR _043_ sky130_fd_sc_hd__and2b_1
XFILLER_0_10_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput19 net19 VGND VGND VPWR VPWR count[6] sky130_fd_sc_hd__buf_1
X_078_ net10 net4 _011_ net16 _028_ VGND VGND VPWR VPWR _003_ sky130_fd_sc_hd__a221o_1
XFILLER_0_2_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_11_Right_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_094_ net12 net19 VGND VGND VPWR VPWR _042_ sky130_fd_sc_hd__and2b_1
XTAP_TAPCELL_ROW_6_33 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_077_ _024_ _026_ _027_ VGND VGND VPWR VPWR _028_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_7_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_4_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_093_ _012_ _039_ _040_ _041_ VGND VGND VPWR VPWR _005_ sky130_fd_sc_hd__a31o_1
XFILLER_0_5_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_3_Left_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput1 data[0] VGND VGND VPWR VPWR net1 sky130_fd_sc_hd__clkbuf_1
X_076_ _024_ _026_ _012_ VGND VGND VPWR VPWR _027_ sky130_fd_sc_hd__o21ai_1
XPHY_EDGE_ROW_9_Right_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_059_ net10 _009_ _011_ _008_ VGND VGND VPWR VPWR _013_ sky130_fd_sc_hd__a22o_1
XFILLER_0_5_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_092_ net10 net6 _011_ net18 VGND VGND VPWR VPWR _041_ sky130_fd_sc_hd__a22o_1
Xinput2 data[1] VGND VGND VPWR VPWR net2 sky130_fd_sc_hd__clkbuf_1
X_075_ net12 _010_ _022_ VGND VGND VPWR VPWR _026_ sky130_fd_sc_hd__o21ai_1
X_058_ net10 net9 VGND VGND VPWR VPWR _012_ sky130_fd_sc_hd__and2b_2
XTAP_TAPCELL_ROW_0_26 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_091_ _037_ _038_ VGND VGND VPWR VPWR _040_ sky130_fd_sc_hd__or2_1
Xinput3 data[2] VGND VGND VPWR VPWR net3 sky130_fd_sc_hd__clkbuf_1
X_074_ _024_ VGND VGND VPWR VPWR _025_ sky130_fd_sc_hd__inv_2
X_057_ net10 net9 VGND VGND VPWR VPWR _011_ sky130_fd_sc_hd__nor2_2
XPHY_EDGE_ROW_0_Right_0 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_12_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_109_ clknet_1_0__leaf_clk _001_ net11 VGND VGND VPWR VPWR net14 sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_0_27 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_9_36 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_090_ _037_ _038_ VGND VGND VPWR VPWR _039_ sky130_fd_sc_hd__nand2_1
Xinput4 data[3] VGND VGND VPWR VPWR net4 sky130_fd_sc_hd__clkbuf_1
X_073_ net12 net16 VGND VGND VPWR VPWR _024_ sky130_fd_sc_hd__xnor2_1
X_056_ net15 VGND VGND VPWR VPWR _010_ sky130_fd_sc_hd__inv_2
X_108_ clknet_1_0__leaf_clk _000_ net11 VGND VGND VPWR VPWR net13 sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_10_37 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput5 data[4] VGND VGND VPWR VPWR net5 sky130_fd_sc_hd__clkbuf_1
X_072_ _012_ _021_ _022_ _023_ VGND VGND VPWR VPWR _002_ sky130_fd_sc_hd__a31o_1
XPHY_EDGE_ROW_10_Left_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_055_ net1 VGND VGND VPWR VPWR _009_ sky130_fd_sc_hd__inv_2
X_107_ _012_ _052_ _053_ VGND VGND VPWR VPWR _007_ sky130_fd_sc_hd__a21o_1
XFILLER_0_11_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput6 data[5] VGND VGND VPWR VPWR net6 sky130_fd_sc_hd__clkbuf_1
X_071_ net10 net3 _011_ net15 VGND VGND VPWR VPWR _023_ sky130_fd_sc_hd__a22o_1
XFILLER_0_2_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_106_ net10 net8 _011_ net20 VGND VGND VPWR VPWR _053_ sky130_fd_sc_hd__a22o_1
X_054_ net13 VGND VGND VPWR VPWR _008_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_4_Right_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput7 data[6] VGND VGND VPWR VPWR net7 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_11_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_070_ _019_ _020_ VGND VGND VPWR VPWR _022_ sky130_fd_sc_hd__or2_1
Xinput10 preload VGND VGND VPWR VPWR net10 sky130_fd_sc_hd__buf_2
X_105_ _050_ _051_ VGND VGND VPWR VPWR _052_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_11_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput8 data[7] VGND VGND VPWR VPWR net8 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_2_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_104_ net12 net20 VGND VGND VPWR VPWR _051_ sky130_fd_sc_hd__xnor2_1
Xinput11 resetn VGND VGND VPWR VPWR net11 sky130_fd_sc_hd__buf_2
Xclkbuf_1_0__f_clk clknet_0_clk VGND VGND VPWR VPWR clknet_1_0__leaf_clk sky130_fd_sc_hd__clkbuf_16
Xinput9 enable VGND VGND VPWR VPWR net9 sky130_fd_sc_hd__buf_1
XPHY_EDGE_ROW_2_Left_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_10_Right_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput12 up_down VGND VGND VPWR VPWR net12 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_2_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_103_ _044_ _046_ _042_ VGND VGND VPWR VPWR _050_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_4_31 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_8_Right_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_102_ _012_ _047_ _048_ _049_ VGND VGND VPWR VPWR _006_ sky130_fd_sc_hd__a31o_1
XFILLER_0_8_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_101_ net10 net7 _011_ net19 VGND VGND VPWR VPWR _049_ sky130_fd_sc_hd__a22o_1
X_100_ _044_ _046_ VGND VGND VPWR VPWR _048_ sky130_fd_sc_hd__or2_1
XPHY_EDGE_ROW_6_Left_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_9_Left_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_8_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_2_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_8_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_7_34 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_61 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_0_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_5_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_3_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_089_ _030_ _033_ _031_ VGND VGND VPWR VPWR _038_ sky130_fd_sc_hd__a21o_1
XFILLER_0_9_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_1_1__f_clk clknet_0_clk VGND VGND VPWR VPWR clknet_1_1__leaf_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_0_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_3_Right_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_6_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_088_ net12 net18 VGND VGND VPWR VPWR _037_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_3_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_12_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_087_ _012_ _034_ _035_ _036_ VGND VGND VPWR VPWR _004_ sky130_fd_sc_hd__a31o_1
XFILLER_0_9_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_1_28 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_086_ net10 net5 _011_ net17 VGND VGND VPWR VPWR _036_ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_1_Left_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_3_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_069_ _019_ _020_ VGND VGND VPWR VPWR _021_ sky130_fd_sc_hd__nand2_1
XPHY_EDGE_ROW_7_Right_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_12_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_11_38 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_085_ _030_ _033_ VGND VGND VPWR VPWR _035_ sky130_fd_sc_hd__nand2_1
XFILLER_0_0_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_068_ net12 net15 VGND VGND VPWR VPWR _020_ sky130_fd_sc_hd__xor2_1
XFILLER_0_12_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_3_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_067_ _008_ _015_ _014_ VGND VGND VPWR VPWR _019_ sky130_fd_sc_hd__o21a_1
X_084_ _030_ _033_ VGND VGND VPWR VPWR _034_ sky130_fd_sc_hd__or2_1
XFILLER_0_12_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_12_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_5_Left_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_083_ _031_ _032_ VGND VGND VPWR VPWR _033_ sky130_fd_sc_hd__nor2_1
XFILLER_0_9_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_8_Left_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_066_ _016_ _017_ _018_ VGND VGND VPWR VPWR _001_ sky130_fd_sc_hd__a21o_1
XFILLER_0_6_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_12_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_12_40 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_065_ net10 net2 _011_ net14 VGND VGND VPWR VPWR _018_ sky130_fd_sc_hd__a22o_1
X_082_ net17 net12 VGND VGND VPWR VPWR _032_ sky130_fd_sc_hd__and2b_1
XFILLER_0_9_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_081_ net12 net17 VGND VGND VPWR VPWR _031_ sky130_fd_sc_hd__and2b_1
XFILLER_0_0_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_064_ _008_ _015_ _012_ VGND VGND VPWR VPWR _017_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_5_32 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_2_Right_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_12_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_2_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_0_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_063_ _008_ _015_ VGND VGND VPWR VPWR _016_ sky130_fd_sc_hd__nand2_1
X_080_ _019_ _020_ _025_ _029_ VGND VGND VPWR VPWR _030_ sky130_fd_sc_hd__o31ai_2
XFILLER_0_10_62 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_115_ clknet_1_1__leaf_clk _007_ net11 VGND VGND VPWR VPWR net20 sky130_fd_sc_hd__dfrtp_1
.ends

