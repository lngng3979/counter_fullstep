VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO counter
  CLASS BLOCK ;
  FOREIGN counter ;
  ORIGIN 0.000 0.000 ;
  SIZE 48.375 BY 59.095 ;
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 24.340 10.640 25.940 46.480 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 46.480 ;
    END
  END VPWR
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 20.440 4.000 21.040 ;
    END
  END clk
  PIN count[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met3 ;
        RECT 44.375 13.640 48.375 14.240 ;
    END
  END count[0]
  PIN count[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 22.630 0.000 22.910 4.000 ;
    END
  END count[1]
  PIN count[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met3 ;
        RECT 0.000 17.040 4.000 17.640 ;
    END
  END count[2]
  PIN count[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met3 ;
        RECT 0.000 27.240 4.000 27.840 ;
    END
  END count[3]
  PIN count[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met3 ;
        RECT 44.375 30.640 48.375 31.240 ;
    END
  END count[4]
  PIN count[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met3 ;
        RECT 44.375 37.440 48.375 38.040 ;
    END
  END count[5]
  PIN count[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 22.630 55.095 22.910 59.095 ;
    END
  END count[6]
  PIN count[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met3 ;
        RECT 0.000 40.840 4.000 41.440 ;
    END
  END count[7]
  PIN data[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 32.290 0.000 32.570 4.000 ;
    END
  END data[0]
  PIN data[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 25.850 0.000 26.130 4.000 ;
    END
  END data[1]
  PIN data[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 16.190 0.000 16.470 4.000 ;
    END
  END data[2]
  PIN data[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 30.640 4.000 31.240 ;
    END
  END data[3]
  PIN data[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 44.375 23.840 48.375 24.440 ;
    END
  END data[4]
  PIN data[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 44.375 34.040 48.375 34.640 ;
    END
  END data[5]
  PIN data[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 25.850 55.095 26.130 59.095 ;
    END
  END data[6]
  PIN data[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 37.440 4.000 38.040 ;
    END
  END data[7]
  PIN enable
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 44.375 27.240 48.375 27.840 ;
    END
  END enable
  PIN preload
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 23.840 4.000 24.440 ;
    END
  END preload
  PIN resetn
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 44.375 17.040 48.375 17.640 ;
    END
  END resetn
  PIN up_down
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 34.040 4.000 34.640 ;
    END
  END up_down
  OBS
      LAYER nwell ;
        RECT 5.330 10.795 42.970 46.430 ;
      LAYER li1 ;
        RECT 5.520 10.795 42.780 46.325 ;
      LAYER met1 ;
        RECT 4.210 10.240 42.780 46.480 ;
      LAYER met2 ;
        RECT 4.230 54.815 22.350 55.095 ;
        RECT 23.190 54.815 25.570 55.095 ;
        RECT 26.410 54.815 41.310 55.095 ;
        RECT 4.230 4.280 41.310 54.815 ;
        RECT 4.230 4.000 15.910 4.280 ;
        RECT 16.750 4.000 22.350 4.280 ;
        RECT 23.190 4.000 25.570 4.280 ;
        RECT 26.410 4.000 32.010 4.280 ;
        RECT 32.850 4.000 41.310 4.280 ;
      LAYER met3 ;
        RECT 3.990 41.840 44.375 46.405 ;
        RECT 4.400 40.440 44.375 41.840 ;
        RECT 3.990 38.440 44.375 40.440 ;
        RECT 4.400 37.040 43.975 38.440 ;
        RECT 3.990 35.040 44.375 37.040 ;
        RECT 4.400 33.640 43.975 35.040 ;
        RECT 3.990 31.640 44.375 33.640 ;
        RECT 4.400 30.240 43.975 31.640 ;
        RECT 3.990 28.240 44.375 30.240 ;
        RECT 4.400 26.840 43.975 28.240 ;
        RECT 3.990 24.840 44.375 26.840 ;
        RECT 4.400 23.440 43.975 24.840 ;
        RECT 3.990 21.440 44.375 23.440 ;
        RECT 4.400 20.040 44.375 21.440 ;
        RECT 3.990 18.040 44.375 20.040 ;
        RECT 4.400 16.640 43.975 18.040 ;
        RECT 3.990 14.640 44.375 16.640 ;
        RECT 3.990 13.240 43.975 14.640 ;
        RECT 3.990 10.715 44.375 13.240 ;
  END
END counter
END LIBRARY

